//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::util::ILocale;

namespace ccm {
namespace io {

/**
 * @Involve interfade ccm::io::IWriter;
 * @Involve interface ccm::core::IAppendable;
 * @Involve interface ccm::io::ICloseable;
 * @Involve interface ccm::io::IFlushable;
 * @involve interface ccm::core::IAutoCloseable
 */
[
    uuid(680fba48-d41b-4a09-9b10-7077eada7b89),
    version(0.1.0)
]
interface IPrintWriter
{
    CheckError(
        [out] Boolean* hasErrors);

    Format(
        [in] String format,
        [in] Array<IInterface*>* args);

    Format(
        [in] ILocale* l,
        [in] String format,
        [in] Array<IInterface*>* args);

    Print(
        [in] Boolean b);

    PrintChar(
        [in] Char c);

    Print(
        [in] Integer i);

    Print(
        [in] Long l);

    Print(
        [in] Float f);

    Print(
        [in] Double d);

    Print(
        [in] Array<Char> s);

    Print(
        [in] String s);

    Print(
        [in] IInterface* obj);

    Printf(
        [in] String format,
        [in] Array<IInterface*>* args);

    Printf(
        [in] ILocale* l,
        [in] String format,
        [in] Array<IInterface*>* args);

    Println();

    Println(
        [in] Boolean b);

    PrintCharln(
        [in] Char c);

    Println(
        [in] Integer i);

    Println(
        [in] Long l);

    Println(
        [in] Float f);

    Println(
        [in] Double x);

    Println(
        [in] Array<Char> s);

    Println(
        [in] String s);

    Println(
        [in] IInterface* obj);
}

}
}
