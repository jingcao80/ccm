//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "util/IArrayList.cdl"
include "util/ICollection.cdl"
include "util/IDictionary.cdl"
include "util/IEnumeration.cdl"
include "util/IHashtable.cdl"
include "util/IIterator.cdl"
include "util/IList.cdl"
include "util/IListIterator.cdl"
include "util/IMap.cdl"
include "util/IRandomAccess.cdl"
include "util/ISet.cdl"
include "util/regex/Exceptions.cdl"
include "util/regex/IMatcher.cdl"
include "util/regex/IMatchResult.cdl"
include "util/regex/IPattern.cdl"

interface ccm::core::ICloneable;
interface ccm::core::IIterable;
interface ccm::io::ISerializable;

namespace ccm {
namespace util {

[
    uuid(7dbd4e0a-4bf2-4ccb-a4e9-bfe232b40ba4),
    version(0.1.0)
]
coclass CArrayList
{
    Constructor();

    interface IArrayList;
    interface IList;
    interface ICollection;
    interface IRandomAccess;
    interface IIterable;
    interface ICloneable;
    interface ISerializable;
}

namespace regex {

[
    uuid(698f1b9a-dd5e-4ae4-924c-c1addd038571),
    version(0.1.0)
]
coclass CPatternFactory
{
    interface IPatternFactory;
}

}
}
}
