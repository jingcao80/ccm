//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace core {

[
    uuid(2108de07-543c-4cc5-9a59-d25121b4568e),
    version(0.1.0)
]
interface IInteger
{
    /**
     * A constant holding the minimum value an {@code int} can
     * have, -2<sup>31</sup>.
     */
    const Integer MIN_VALUE = 0x80000000;

    /**
     * A constant holding the maximum value an {@code int} can
     * have, 2<sup>31</sup>-1.
     */
    const Integer MAX_VALUE = 0x7fffffff;

    ByteValue(
        [out] Byte* value);

    CompareTo(
        [in] IInterface* other,
        [out] Integer* result);

    DoubleValue(
        [out] Double* value);

    FloatValue(
        [out] Float* value);

    GetValue(
        [out] Integer* value);

    IntValue(
        [out] Integer* value);

    LongValue(
        [out] Long* value);

    ShortValue(
        [out] Short* value);
}

}
}
