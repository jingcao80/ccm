//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace io {

const Integer E_IO_EXCEPTION = 0x80010200;
const Integer E_IO_SYNC_FAILED_EXCEPTION = 0x80010201;
const Integer E_FILE_NOT_FOUND_EXCEPTION = 0x80010202;
const Integer E_USE_MANUAL_SKIP_EXCEPTION = 0x80010203;

}
}