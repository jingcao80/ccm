//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "core/Errors.cdl"
include "core/Exceptions.cdl"
include "core/IAppendable.cdl"
include "core/IArray.cdl"
include "core/IBoolean.cdl"
include "core/IByte.cdl"
include "core/IChar.cdl"
include "core/ICharSequence.cdl"
include "core/ICloneable.cdl"
include "core/IComparable.cdl"
include "core/IDouble.cdl"
include "core/IFloat.cdl"
include "core/IInteger.cdl"
include "core/IIterable.cdl"
include "core/ILong.cdl"
include "core/INumber.cdl"
include "core/IRunnable.cdl"
include "core/IShort.cdl"
include "core/IStackTraceElement.cdl"
include "core/IString.cdl"
include "core/IStringBuffer.cdl"
include "core/IStringBuilder.cdl"
include "core/ISynchronize.cdl"
include "core/IThread.cdl"
include "core/IThreadGroup.cdl"

namespace ccm {
namespace core {

[
    uuid(bc5be123-34ab-4373-ab98-31c3e3c68b1b),
    version(0.1.0)
]
coclass CArray
{
    Constructor(
        [in] InterfaceID elemId,
        [in] Long size);

    interface IArray;
}

[
    uuid(339a8069-7448-4d12-9c50-d45497fb245b),
    version(0.1.0)
]
coclass CThread
{
    Constructor();

    Constructor(
        [in] IThreadGroup* group,
        [in] String name,
        [in] Integer priority,
        [in] Boolean daemon);

    // @hide
    Constructor(
        [in] HANDLE peer);

    interface IRunnable;
    interface IThread;
}

[
    uuid(730c7375-05c3-4b86-933c-ab2808164280),
    version(0.1.0)
]
coclass CThreadGroup
{
    // @hide
    Constructor();

    Constructor(
        [in] String name);

    Constructor(
        [in] IThreadGroup* parent,
        [in] String name);

    interface IThreadGroup;
}

}
}
