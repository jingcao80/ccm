//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace core {

/*
 * @Involve interface como::core::INumber
 * @Involve interface como::core::IComparable
 * @Involve interface como::io::ISerializable
 */
[
    uuid(b0acf41b-e045-461e-88a4-64c1486ac78a),
    version(0.1.0)
]
interface ILong
{
    /**
     * A constant holding the minimum value a {@code long} can
     * have, -2<sup>63</sup>.
     */
    const Long MIN_VALUE = 0x8000000000000000ll;

    /**
     * A constant holding the maximum value a {@code long} can
     * have, 2<sup>63</sup>-1.
     */
    const Long MAX_VALUE = 0x7fffffffffffffffll;

    const Integer SIZE = 64;

    ByteValue(
        [out] Byte& value);

    CompareTo(
        [in] IInterface* other,
        [out] Integer& result);

    DoubleValue(
        [out] Double& value);

    FloatValue(
        [out] Float& value);

    GetValue(
        [out] Long& value);

    IntegerValue(
        [out] Integer& value);

    LongValue(
        [out] Long& value);

    ShortValue(
        [out] Short& value);
}

}
}
