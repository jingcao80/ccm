//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::util::ICollection;

namespace como {
namespace util {

/*
 * @Involve interface como::util::IList;
 * @Involve interface como::util::ICollection;
 * @Involve interface como::core::IIterable;
 * @Involve interface como::util::IDeque;
 * @Involve interface como::util::IQueue;
 */
[
    uuid(116514aa-3d9b-480a-a3f1-77b8cfab8ae2),
    version(0.1.0)
]
interface ILinkedList
{
    Add(
        [in] IInterface* e,
        [out] Boolean* changed = nullptr);

    Add(
        [in] Integer index,
        [in] IInterface* obj);

    AddAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    AddAll(
        [in] Integer index,
        [in] ICollection* c,
        [out] Boolean* result = nullptr);

    AddFirst(
        [in] IInterface* e);

    AddLast(
        [in] IInterface* e);

    Clear();

    Contains(
        [in] IInterface* obj,
        [out] Boolean& result);

    Element(
        [out] IInterface&& e);

    Get(
        [in] Integer index,
        [out] IInterface** obj);

    GetFirst(
        [out] IInterface** e);

    GetIterator(
        [out] IIterator&& it);

    GetLast(
        [out] IInterface** e);

    GetListIterator(
        [in] Integer index,
        [out] IListIterator** it);

    GetSize(
        [out] Integer& size);

    IndexOf(
        [in] IInterface* obj,
        [out] Integer* index);

    LastIndexOf(
        [in] IInterface* obj,
        [out] Integer* index);

    Offer(
        [in] IInterface* e,
        [out] Boolean* changed = nullptr);

    OfferFirst(
        [in] IInterface* e,
        [out] Boolean* changed = nullptr);

    OfferLast(
        [in] IInterface* e,
        [out] Boolean* changed = nullptr);

    Peek(
        [out] IInterface&& e);

    PeekFirst(
        [out] IInterface** e);

    PeekLast(
        [out] IInterface** e);

    Poll(
        [out] IInterface** e);

    PollFirst(
        [out] IInterface** e);

    PollLast(
        [out] IInterface** e);

    Pop(
        [out] IInterface** e);

    Push(
        [in] IInterface* e);

    Remove(
        [out] IInterface** e = nullptr);

    Remove(
        [in] IInterface* obj,
        [out] Boolean* result = nullptr);

    Remove(
        [in] Integer index,
        [out] IInterface** obj = nullptr);

    RemoveFirst(
        [out] IInterface** e = nullptr);

    RemoveFirstOccurrence(
        [in] IInterface* e,
        [out] Boolean* changed = nullptr);

    RemoveLast(
        [out] IInterface** e = nullptr);

    RemoveLastOccurrence(
        [in] IInterface* e,
        [out] Boolean* changed = nullptr);

    Set(
        [in] Integer index,
        [in] IInterface* obj,
        [out] IInterface** prevObj = nullptr);
}

}
}
