//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {

[
    uuid(6a87e3db-c2aa-470c-9638-4a2d31dfdd35),
    version(0.1.0)
]
interface IDate
{
    After(
        [in] IDate* when,
        [out] Boolean* after);

    Before(
        [in] IDate* when,
        [out] Boolean* before);

    GetDate(
        [out] Integer* date);

    GetDay(
        [out] Integer* day);

    GetHours(
        [out] Integer* hours);

    GetMinutes(
        [out] Integer* minutes);

    GetMonth(
        [out] Integer* month);

    GetSeconds(
        [out] Integer* seconds);

    GetTime(
        [out] Long* time);

    GetTimezoneOffset(
        [out] Integer* tzOffset);

    GetYear(
        [out] Integer* year);

    SetDate(
        [in] Integer date);

    SetHours(
        [in] Integer hours);

    SetMinutes(
        [in] Integer minutes);

    SetMonth(
        [in] Integer month);

    SetSeconds(
        [in] Integer seconds);

    SetTime(
        [in] Long time);

    SetYear(
        [in] Integer year);

    ToGMTString(
        [out] String* str);

    ToLocaleString(
        [out] String* str);
}

}
}
