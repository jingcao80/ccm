//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {

/*
 * @Involve interface como::util::IEnumeration
 */
[
    uuid(8283c934-d3ce-4a7b-ad50-a97f757ce121),
    version(0.1.0)
]
interface IStringTokenizer
{
    CountTokens(
        [out] Integer& number);

    HasMoreElements(
        [out] Boolean& hasMore);

    HasMoreTokens(
        [out] Boolean& hasMore);

    NextElement(
        [out] IInterface&& element);

    NextToken(
        [out] String& token);

    NextToken(
        [in] String delim,
        [out] String& token);
}

}
}
