//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::core::IStringBuffer;
interface como::text::IFieldPosition;

namespace como {
namespace text {

/*
 * @Involve interface como::text::INumberFormat;
 * @Involve interface como::text::IFormat;
 * @Involve interface como::io::ISerializable;
 * @Involve interface como::core::ICloneable;
 */
[
    uuid(54f82f1f-4aaf-45b6-891d-77083bff1058),
    version(0.1.0)
]
interface IChoiceFormat
{
    ApplyPattern(
        [in] String newPattern);

    Format(
        [in] Long number,
        [out] IStringBuffer* toAppendTo,
        [in] IFieldPosition* status);

    Format(
        [in] Double number,
        [out] IStringBuffer* toAppendTo,
        [in] IFieldPosition* status);

    GetFormats(
        [out, callee] Array<String>* formats);

    GetLimits(
        [out, callee] Array<Double>* limits);

    SetChoices(
        [in] Array<Double> limits,
        [in] Array<String> formats);

    ToPattern(
        [out] String& pattern);
}

}
}
