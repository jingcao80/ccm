//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace core {

[
    uuid(7ddf21a8-3891-484e-a23b-2ad9cedabf17),
    version(0.1.0)
]
interface ISynchronize
{
    Lock();

    Unlock();

    Notify();

    NotifyAll();

    Wait();

    Wait(
        [in] Long millis);

    Wait(
        [in] Long millis,
        [in] Integer nanos);
}

}
}
