//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace io {

[
    uuid(23485c78-6782-4d5f-8d30-55cf6a6e5dde),
    version(0.1.0)
]
interface IDoubleBuffer
{
    AsReadOnlyBuffer(
        [out] IDoubleBuffer&& buffer);

    Compact();

    Duplicate(
        [out] IDoubleBuffer&& buffer);

    Get(
        [out] Double& d);

    Get(
        [in] Integer index,
        [out] Double& d);

    Get(
        [out] Array<Double>& dst);

    Get(
        [out] Array<Double>& dst,
        [in] Integer offset,
        [in] Integer length);

    GetOrder(
        [out] IByteOrder&& bo);

    HasArray(
        [out] Boolean& result);

    Put(
        [in] Double d);

    Put(
        [in] Integer index,
        [in] Double d);

    Put(
        [in] Array<Double> src);

    Put(
        [in] Array<Double> src,
        [in] Integer offset,
        [in] Integer length);

    Put(
        [in] IDoubleBuffer* src);

    Slice(
        [out] IDoubleBuffer&& buffer);
}

}
}
