//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ccm/io/Exceptions.cdl"
include "ccm/io/IBuffer.cdl"
include "ccm/io/IBufferedWriter.cdl"
include "ccm/io/IByteArrayOutputStream.cdl"
include "ccm/io/IByteBuffer.cdl"
include "ccm/io/IByteOrder.cdl"
include "ccm/io/ICharBuffer.cdl"
include "ccm/io/ICloseable.cdl"
include "ccm/io/IDoubleBuffer.cdl"
include "ccm/io/IFile.cdl"
include "ccm/io/IFileDescriptor.cdl"
include "ccm/io/IFileFilter.cdl"
include "ccm/io/IFileInputStream.cdl"
include "ccm/io/IFileOutputStream.cdl"
include "ccm/io/IFilenameFilter.cdl"
include "ccm/io/IFloatBuffer.cdl"
include "ccm/io/IFlushable.cdl"
include "ccm/io/IInputStream.cdl"
include "ccm/io/IIntegerBuffer.cdl"
include "ccm/io/IInterruptible.cdl"
include "ccm/io/ILongBuffer.cdl"
include "ccm/io/IMappedByteBuffer.cdl"
include "ccm/io/IOutputStream.cdl"
include "ccm/io/IOutputStreamWriter.cdl"
include "ccm/io/IPrintStream.cdl"
include "ccm/io/IPrintWriter.cdl"
include "ccm/io/IReader.cdl"
include "ccm/io/ISerializable.cdl"
include "ccm/io/IShortBuffer.cdl"
include "ccm/io/IStringWriter.cdl"
include "ccm/io/IWriter.cdl"
include "ccm/io/channels/IDirectBuffer.cdl"
include "ccm/io/channels/IFileChannel.cdl"
include "ccm/io/charset/ICharset.cdl"
include "ccm/io/charset/ICharsetEncoder.cdl"
include "ccm/io/charset/IStreamEncoder.cdl"

interface ccm::core::IAppendable;
interface ccm::core::IAutoCloseable;
interface ccm::core::IComparable;
interface ccm::io::channels::IDirectBuffer;
interface ccm::io::charset::ICharset;
interface ccm::io::charset::ICharsetEncoder;
interface ccm::net::IURI;

namespace ccm {
namespace io {

[
    uuid(cf7b3ffb-46ce-44fc-9057-d8ec03c820b7),
    version(0.1.0)
]
coclass CBufferedWriter
{
    Constructor(
        [in] IWriter* outW);

    Constructor(
        [in] IWriter* outW,
        [in] Integer sz);

    interface IBufferedWriter;
    interface IWriter;
    interface IAppendable;
    interface ICloseable;
    interface IFlushable;
    interface IAutoCloseable;
}

[
    uuid(69455e4d-56b1-43b1-98b1-e4907e332a4f),
    version(0.1.0)
]
coclass CByteArrayOutputStream
{
    Constructor();

    Constructor(
        [in] Integer size);

    interface IByteArrayOutputStream;
    interface IOutputStream;
    interface IFlushable;
    interface ICloseable;
    interface IAutoCloseable;
}

[
    uuid(160997fd-1165-46dd-a47a-8a000bcd1916),
    version(0.1.0)
]
coclass CDirectByteBuffer
{
    Constructor(
        [in] Integer cap,
        [in] HANDLE address,
        [in] IFileDescriptor* fd,
        [in] Boolean isReadOnly);

    interface IDirectBuffer;
    interface IMappedByteBuffer;
    interface IByteBuffer;
    interface IBuffer;
    interface IComparable;
}

[
    uuid(0d9c5571-7eaa-44e1-815f-c6af421c780d),
    version(0.1.0)
]
coclass CFile
{
    Constructor(
        [in] String pathname);

    Constructor(
        [in] String parent,
        [in] String child);

    Constructor(
        [in] IFile* parent,
        [in] String child);

    Constructor(
        [in] IURI* uri);

    // @hide
    Constructor(
        [in] String pathname,
        [in] Integer prefixLength);

    // @hide
    Constructor(
        [in] String child,
        [in] IFile* parent);

    interface IFile;
}

[
    uuid(3e291dd3-0c31-4526-8ef9-fe61bc1e508e),
    version(0.1.0)
]
coclass CFileDescriptor
{
    Constructor();

    Constructor(
        [in] Integer descriptor);

    interface IFileDescriptor;
}

[
    uuid(28063bc3-48b2-43f4-b159-c4c65475b844),
    version(0.1.0)
]
coclass CFileInputStream
{
    Constructor(
        [in] String name);

    Constructor(
        [in] IFile* file);

    Constructor(
        [in] IFileDescriptor* fdObj);

    Constructor(
        [in] IFileDescriptor* fdObj,
        [in] Boolean isFdOwner);

    interface IFileInputStream;
    interface IInputStream;
    interface ICloseable;
    interface IAutoCloseable;
}

[
    uuid(6d5f9b98-ce5c-4e30-a5ca-c0c74e0dc8fd),
    version(0.1.0)
]
coclass CFileOutputStream
{
    Constructor(
        [in] String name);

    Constructor(
        [in] String name,
        [in] Boolean append);

    Constructor(
        [in] IFile* file);

    Constructor(
        [in] IFile* file,
        [in] Boolean append);

    Constructor(
        [in] IFileDescriptor* fdObj);

    Constructor(
        [in] IFileDescriptor* fdObj,
        [in] Boolean isFdOwner);

    interface IFileOutputStream;
    interface IOutputStream;
    interface IFlushable;
    interface ICloseable;
    interface IAutoCloseable;
}

[
    uuid(3f1442a5-ce76-40b3-8889-c9431c810c1d),
    version(0.1.0)
]
coclass COutputStreamWriter
{
    Constructor(
        [in] IOutputStream* outstream,
        [in] String charsetName);

    Constructor(
        [in] IOutputStream* outstream);

    Constructor(
        [in] IOutputStream* outstream,
        [in] ICharset* cs);

    Constructor(
        [in] IOutputStream* outstream,
        [in] ICharsetEncoder* enc);

    interface IOutputStreamWriter;
    interface IWriter;
    interface IAppendable;
    interface ICloseable;
    interface IFlushable;
    interface IAutoCloseable;
}

[
    uuid(5de87670-f240-43cd-b06d-a758b4914e76),
    version(0.1.0)
]
coclass CPrintWriter
{
    Constructor(
        [in] IWriter* outstream);

    Constructor(
        [in] IWriter* outstream,
        [in] Boolean autoFlush);

    Constructor(
        [in] IOutputStream* outstream);

    Constructor(
        [in] IOutputStream* outstream,
        [in] Boolean autoFlush);

    Constructor(
        [in] String fileName);

    Constructor(
        [in] String fileName,
        [in] String csn);

    Constructor(
        [in] IFile* file);

    Constructor(
        [in] IFile* file,
        [in] String csn);

    interface IPrintWriter;
}

[
    uuid(2a886435-1ec8-4311-be20-03cff45b0dc8),
    version(0.1.0)
]
coclass CStringWriter
{
    Constructor();

    Constructor(
        [in] Integer initialSize);

    interface IStringWriter;
    interface IWriter;
    interface IAppendable;
    interface ICloseable;
    interface IFlushable;
    interface IAutoCloseable;
}

}
}
