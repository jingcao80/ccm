//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::util::ICurrency;

namespace como {
namespace text {

/*
 * @Involve interface como::io::ISerializable
 * @Involve interface como::core::ICloneable
 */
[
    uuid(e7a8ca7c-5f0b-4d11-b50e-25d3593720d8),
    version(0.1.0)
]
interface IDecimalFormatSymbols
{
    GetCurrency(
        [out] ICurrency&& currency);

    GetCurrencySymbol(
        [out] String& currency);

    GetDecimalSeparator(
        [out] Char& decimalSeparator);

    GetDigit(
        [out] Char& digit);

    GetExponentSeparator(
        [out] String& exponentSeparator);

    GetGroupingSeparator(
        [out] Char& groupingSeparator);

    GetInfinity(
        [out] String& infinity);

    GetInternationalCurrencySymbol(
        [out] String& currency);

    GetMinusSign(
        [out] Char& minusSign);

    GetMinusSignString(
        [out] String& minusSignStr);

    GetMonetaryDecimalSeparator(
        [out] Char& monetarySeparator);

    GetNaN(
        [out] String& naN);

    GetPatternSeparator(
        [out] Char& patternSeparator);

    GetPercent(
        [out] Char& percent);

    GetPercentString(
        [out] String& percentStr);

    GetPerMill(
        [out] Char& perMill);

    GetZeroDigit(
        [out] Char& zeroDigit);

    SetCurrency(
        [in] ICurrency* currency);

    SetCurrencySymbol(
        [in] String currency);

    SetDecimalSeparator(
        [in] Char decimalSeparator);

    SetDigit(
        [in] Char digit);

    SetExponentSeparator(
        [in] String exp);

    SetGroupingSeparator(
        [in] Char groupingSeparator);

    SetInfinity(
        [in] String infinity);

    SetInternationalCurrencySymbol(
        [in] String currency);

    SetMinusSign(
        [in] Char minusSign);

    SetMonetaryDecimalSeparator(
        [in] Char sep);

    SetNaN(
        [in] String naN);

    SetPatternSeparator(
        [in] Char patternSeparator);

    SetPercent(
        [in] Char percent);

    SetPerMill(
        [in] Char perMill);

    SetZeroDigit(
        [in] Char zeroDigit);
}

}
}
