//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface libcore::io::IBufferIterator;

namespace libcore {
namespace io {

/*
 * @Involve interface como::core::IAutoCloseable;
 */
[
    uuid(c3142383-5fa7-4fe7-a98e-c5e5bf321c58),
    version(0.1.0)
]
interface IMemoryMappedFile
{
    BigEndianIterator(
        [out] IBufferIterator** it);

    IsClosed(
        [out] Boolean* closed);

    LittleEndianIterator(
        [out] IBufferIterator** it);

    GetSize(
        [out] Integer* size);
}

}
}
