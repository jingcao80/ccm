//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ccm/security/IGuard.cdl"
include "ccm/security/IPermission.cdl"
include "ccm/security/IPermissionCollection.cdl"
include "ccm/security/IPrivilegedAction.cdl"

namespace ccm {
namespace security {

namespace action {

[
    uuid(b2412c80-ec7f-46de-a4de-6ade765814da),
    version(0.1.0)
]
coclass CGetPropertyAction
{
    Constructor(
        [in] String theProp);

    Constructor(
        [in] String theProp
        [in] String defaultVal);

    interface IPrivilegedAction;
}

}

}
}
