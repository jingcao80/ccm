//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::io::IFileFilter;
interface como::io::IFilenameFilter;
interface como::net::IURI;
interface como::net::IURL;

namespace como {
namespace io {

/*
 * @Involve interface como::core::IComparable
 * @Involve interface como::io::ISerializable
 */
[
    uuid(64d64034-3b89-4cc0-b446-d20c3a6a0f8f),
    version(0.1.0)
]
interface IFile
{
    CanExecute(
        [out] Boolean* executable);

    CanRead(
        [out] Boolean* readable);

    CanWrite(
        [out] Boolean* writeable);

    CreateNewFile(
        [out] Boolean* succeeded);

    Delete(
        [out] Boolean* succeeded = nullptr);

    DeleteOnExit();

    Exists(
        [out] Boolean* existed);

    GetAbsoluteFile(
        [out] IFile** f);

    GetAbsolutePath(
        [out] String* path);

    GetCanonicalFile(
        [out] IFile** f);

    GetCanonicalPath(
        [out] String* path);

    GetFreeSpace(
        [out] Long* space);

    GetLength(
        [out] Long* len);

    GetName(
        [out] String* name);

    GetParent(
        [out] String* parent);

    GetParentFile(
        [out] IFile** parent);

    GetPath(
        [out] String* path);

    // @hide
    GetPrefixLength(
        [out] Integer* length);

    GetTotalSpace(
        [out] Long* space);

    GetUsableSpace(
        [out] Long* space);

    IsAbsolute(
        [out] Boolean* absolute);

    IsDirectory(
        [out] Boolean* directory);

    IsFile(
        [out] Boolean* file);

    IsHidden(
        [out] Boolean* hidden);

    LastModified(
        [out] Long* time);

    List(
        [out, callee] Array<String>* files);

    List(
        [in] IFilenameFilter* filter,
        [out, callee] Array<String>* files);

    ListFiles(
        [out, callee] Array<IFile*>* files);

    ListFiles(
        [in] IFilenameFilter* filter,
        [out, callee] Array<IFile*>* files);

    ListFiles(
        [in] IFileFilter* filter,
        [out, callee] Array<IFile*>* files);

    Mkdir(
        [out] Boolean* succeeded);

    Mkdirs(
        [out] Boolean* succeeded);

    RenameTo(
        [in] IFile* dest,
        [out] Boolean* succeeded);

    SetExecutable(
        [in] Boolean executable,
        [out] Boolean* succeeded);

    SetExecutable(
        [in] Boolean executable,
        [in] Boolean ownerOnly,
        [out] Boolean* succeeded);

    SetLastModified(
        [in] Long time,
        [out] Boolean* succeeded);

    SetReadOnly(
        [out] Boolean* succeeded);

    SetReadable(
        [in] Boolean readable,
        [out] Boolean* succeeded);

    SetReadable(
        [in] Boolean readable,
        [in] Boolean ownerOnly,
        [out] Boolean* succeeded);

    SetWritable(
        [in] Boolean writable,
        [out] Boolean* succeeded);

    SetWritable(
        [in] Boolean writable,
        [in] Boolean ownerOnly,
        [out] Boolean* succeeded);

    ToURI(
        [out] IURI** id);

    ToURL(
        [out] IURL** locator);
}

}
}
