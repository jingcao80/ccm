//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::IArgumentList;
interface como::IClassLoader;
interface como::IMetaCoclass;
interface como::IMetaConstant;
interface como::IMetaConstructor;
interface como::IMetaEnumeration;
interface como::IMetaEnumerator;
interface como::IMetaInterface;
interface como::IMetaMethod;
interface como::IMetaParameter;
interface como::IMetaType;
interface como::IMetaValue;

namespace como {

enum IOAttribute
{
    UNKNOWN,
    IN,
    OUT,
    IN_OUT,
    OUT_CALLEE
}

[
    uuid(35b4d7ca-b66c-44d3-b4a6-007852953085),
    version(0.1.0)
]
interface IMetaComponent
{
    GetName(
        [out] String& name);

    GetComponentID(
        [out] ComponentID& cid);

    GetCoclassNumber(
        [out] Integer& number);

    GetAllCoclasses(
        [out] Array<IMetaCoclass*>& klasses);

    GetCoclass(
        [in] String fullName,
        [out] IMetaCoclass&& klass);

    GetCoclass(
        [in] CoclassID cid,
        [out] IMetaCoclass&& klass);

    GetInterfaceNumber(
        [out] Integer& number);

    GetAllInterfaces(
        [out] Array<IMetaInterface*>& intfs);

    GetInterface(
        [in] String fullName,
        [out] IMetaInterface&& intf);

    GetInterface(
        [in] InterfaceID iid,
        [out] IMetaInterface&& intf);

    GetEnumerationNumber(
        [out] Integer& number);

    GetAllEnumerations(
        [out] Array<IMetaEnumeration*>& enumns);

    GetEnumeration(
        [in] String fullName,
        [out] IMetaEnumeration&& enumn);

    CanUnload(
        [out] Boolean& unload);

    Unload();
}

[
    uuid(8fdbd639-39be-4e9f-801d-8a3b137d7c1f),
    version(0.1.0)
]
interface IMetaCoclass
{
    GetComponent(
        [out] IMetaComponent&& comp);

    GetName(
        [out] String& name);

    GetNamespace(
        [out] String& ns);

    GetCoclassID(
        [out] CoclassID& cid);

    GetClassLoader(
        [out] IClassLoader&& loader);

    GetConstructorNumber(
        [out] Integer& number);

    GetAllConstructors(
        [out] Array<IMetaConstructor*>& constrs);

    GetConstructor(
        [in] String signature,
        [out] IMetaConstructor&& constr);

    GetInterfaceNumber(
        [out] Integer& number);

    GetAllInterfaces(
        [out] Array<IMetaInterface*>& intfs);

    GetInterface(
        [in] String fullName,
        [out] IMetaInterface&& intf);

    ContainsInterface(
        [in] String fullName,
        [out] Boolean& result);

    GetMethodNumber(
        [out] Integer& number);

    GetAllMethods(
        [out] Array<IMetaMethod*>& methods);

    GetMethod(
        [in] String name,
        [in] String signature,
        [out] IMetaMethod&& method);

    CreateObject(
        [in] InterfaceID iid,
        [out] IInterface&& object);
}

[
    uuid(f23514ea-5b7f-4a16-85da-102decb85d38),
    version(0.1.0)
]
interface IMetaEnumeration
{
    GetComponent(
        [out] IMetaComponent&& comp);

    GetName(
        [out] String& name);

    GetNamespace(
        [out] String& ns);

    GetEnumeratorNumber(
        [out] Integer& number);

    GetAllEnumerators(
        [out] Array<IMetaEnumerator*>& enumrs);

    GetEnumerator(
        [in] String name,
        [out] IMetaEnumerator&& enumr);
}

[
    uuid(f508e549-ba3f-4a6e-ad4b-b8bdd3c3fe73),
    version(0.1.0)
]
interface IMetaEnumerator
{
    GetEnumeration(
        [out] IMetaEnumeration&& enumn);

    GetName(
        [out] String& name);

    GetValue(
        [out] Integer& value);
}

[
    uuid(a9f54826-5903-4910-af5f-9703364663b2),
    version(0.1.0)
]
interface IMetaInterface
{
    GetComponent(
        [out] IMetaComponent&& comp);

    GetName(
        [out] String& name);

    GetNamespace(
        [out] String& ns);

    GetInterfaceID(
        [out] InterfaceID& iid);

    GetBaseInterface(
        [out] IMetaInterface&& baseIntf);

    GetConstantNumber(
        [out] Integer& number);

    GetAllConstants(
        [out] Array<IMetaConstant*>& consts);

    GetConstant(
        [in] String name,
        [out] IMetaConstant&& constt);

    GetConstant(
        [in] Integer index,
        [out] IMetaConstant&& constt);

    GetMethodNumber(
        [out] Integer& number);

    GetAllMethods(
        [out] Array<IMetaMethod*>& methods);

    GetMethod(
        [in] String name,
        [in] String signature,
        [out] IMetaMethod&& method);

    GetMethod(
        [in] Integer index,
        [out] IMetaMethod&& method);
}

[
    uuid(c27054e4-f998-4eac-9a2c-17d05aa6dccd),
    version(0.1.0)
]
interface IMetaConstant
{
    GetName(
        [out] String& name);

    GetType(
        [out] IMetaType&& type);

    GetValue(
        [out] IMetaValue&& value);
}

[
    uuid(684f21a0-6d9f-4784-b641-c74fb71c530a),
    version(0.1.0)
]
interface IMetaMethod
{
    GetInterface(
        [out] IMetaInterface&& intf);

    GetName(
        [out] String& name);

    GetSignature(
        [out] String& signature);

    GetParameterNumber(
        [out] Integer& number);

    GetAllParameters(
        [out] Array<IMetaParameter*>& params);

    GetParameter(
        [in] Integer index,
        [out] IMetaParameter&& param);

    GetParameter(
        [in] String name,
        [out] IMetaParameter&& param);

    HasOutArguments(
        [out] Boolean& outArgs);

    CreateArgumentList(
        [out] IArgumentList&& argList);

    Invoke(
        [in] IInterface* thisObject,
        [in] IArgumentList* argList);
}

[
    uuid(ba7707a3-e2f8-4318-8559-f12940f02b2e),
    version(0.1.0)
]
interface IMetaConstructor : IMetaMethod
{
    GetCoclass(
        [out] IMetaCoclass&& klass);

    IsDefault(
        [out] Boolean& isDefault);

    CreateObject(
        [in] IArgumentList* argList,
        [out] IInterface&& object);
}

[
    uuid(0f1060f0-93ea-4980-96b3-bea869dcf253),
    version(0.1.0)
]
interface IMetaParameter
{
    GetMethod(
        [out] IMetaMethod&& method);

    GetName(
        [out] String& name);

    GetIndex(
        [out] Integer& index);

    GetIOAttribute(
        [out] IOAttribute& attr);

    GetType(
        [out] IMetaType&& type);
}

[
    uuid(c9e137d6-2344-4acb-9a76-4d0a9dea1773),
    version(0.1.0)
]
interface IMetaType
{
    GetName(
        [out] String& name);

    GetTypeKind(
        [out] Integer& kind);

    GetElementType(
        [out] IMetaType&& elemType);

    GetPointerNumber(
        [out] Integer& number);
}

[
    uuid(c0dfe841-80a0-421c-ad0a-be51c9d2a0c9),
    version(0.1.0)
]
interface IMetaValue
{
    GetType(
        [out] IMetaType&& type);

    GetBooleanValue(
        [out] Boolean& value);

    GetCharValue(
        [out] Char& value);

    GetByteValue(
        [out] Byte& value);

    GetShortValue(
        [out] Short& value);

    GetIntegerValue(
        [out] Integer& value);

    GetLongValue(
        [out] Long& value);

    GetFloatValue(
        [out] Float& value);

    GetDoubleValue(
        [out] Double& value);

    GetStringValue(
        [out] String& value);

    GetRadix(
        [out] Integer& radix);
}

[
    uuid(38c359ba-97b3-4b7b-bcf7-cd5f6bbed6e9),
    version(0.1.0)
]
interface IArgumentList
{
    GetInputArgumentOfByte(
        [in] Integer index,
        [out] Byte& value);

    SetInputArgumentOfByte(
        [in] Integer index,
        [in] Byte value);

    GetInputArgumentOfShort(
        [in] Integer index,
        [out] Short& value);

    SetInputArgumentOfShort(
        [in] Integer index,
        [in] Short value);

    GetInputArgumentOfInteger(
        [in] Integer index,
        [out] Integer& value);

    SetInputArgumentOfInteger(
        [in] Integer index,
        [in] Integer value);

    GetInputArgumentOfLong(
        [in] Integer index,
        [out] Long& value);

    SetInputArgumentOfLong(
        [in] Integer index,
        [in] Long value);

    GetInputArgumentOfFloat(
        [in] Integer index,
        [out] Float& value);

    SetInputArgumentOfFloat(
        [in] Integer index,
        [in] Float value);

    GetInputArgumentOfDouble(
        [in] Integer index,
        [out] Double& value);

    SetInputArgumentOfDouble(
        [in] Integer index,
        [in] Double value);

    GetInputArgumentOfChar(
        [in] Integer index,
        [out] Char& value);

    SetInputArgumentOfChar(
        [in] Integer index,
        [in] Char value);

    GetInputArgumentOfBoolean(
        [in] Integer index,
        [out] Boolean& value);

    SetInputArgumentOfBoolean(
        [in] Integer index,
        [in] Boolean value);

    GetInputArgumentOfString(
        [in] Integer index,
        [out] String& value);

    SetInputArgumentOfString(
        [in] Integer index,
        [in] String value);

    GetInputArgumentOfHANDLE(
        [in] Integer index,
        [out] HANDLE& value);

    SetInputArgumentOfHANDLE(
        [in] Integer index,
        [in] HANDLE value);

    GetInputArgumentOfECode(
        [in] Integer index,
        [out] ECode& value);

    SetInputArgumentOfECode(
        [in] Integer index,
        [in] ECode value);

    GetInputArgumentOfCoclassID(
        [in] Integer index,
        [out] CoclassID& value);

    SetInputArgumentOfCoclassID(
        [in] Integer index,
        [in] CoclassID value);

    GetInputArgumentOfComponentID(
        [in] Integer index,
        [out] ComponentID& value);

    SetInputArgumentOfComponentID(
        [in] Integer index,
        [in] ComponentID value);

    GetInputArgumentOfInterfaceID(
        [in] Integer index,
        [out] InterfaceID& value);

    SetInputArgumentOfInterfaceID(
        [in] Integer index,
        [in] InterfaceID value);

    GetInputArgumentOfArray(
        [in] Integer index,
        [out] HANDLE& value);

    SetInputArgumentOfArray(
        [in] Integer index,
        [in] HANDLE value);

    GetInputArgumentOfEnumeration(
        [in] Integer index,
        [out] Integer& value);

    SetInputArgumentOfEnumeration(
        [in] Integer index,
        [in] Integer value);

    GetInputArgumentOfInterface(
        [in] Integer index,
        [out] IInterface&& value);

    SetInputArgumentOfInterface(
        [in] Integer index,
        [in] IInterface* value);

    AssignOutputArgumentOfByte(
        [in] Integer index,
        [in] Byte value);

    SetOutputArgumentOfByte(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfShort(
        [in] Integer index,
        [in] Short value);

    SetOutputArgumentOfShort(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfInteger(
        [in] Integer index,
        [in] Integer value);

    SetOutputArgumentOfInteger(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfLong(
        [in] Integer index,
        [in] Long value);

    SetOutputArgumentOfLong(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfFloat(
        [in] Integer index,
        [in] Float value);

    SetOutputArgumentOfFloat(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfDouble(
        [in] Integer index,
        [in] Double value);

    SetOutputArgumentOfDouble(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfChar(
        [in] Integer index,
        [in] Char value);

    SetOutputArgumentOfChar(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfBoolean(
        [in] Integer index,
        [in] Boolean value);

    SetOutputArgumentOfBoolean(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfString(
        [in] Integer index,
        [in] String value);

    SetOutputArgumentOfString(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfHANDLE(
        [in] Integer index,
        [in] HANDLE value);

    SetOutputArgumentOfHANDLE(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfECode(
        [in] Integer index,
        [in] ECode value);

    SetOutputArgumentOfECode(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfCoclassID(
        [in] Integer index,
        [in] CoclassID value);

    SetOutputArgumentOfCoclassID(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfComponentID(
        [in] Integer index,
        [in] ComponentID value);

    SetOutputArgumentOfComponentID(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfInterfaceID(
        [in] Integer index,
        [in] InterfaceID value);

    SetOutputArgumentOfInterfaceID(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfArray(
        [in] Integer index,
        [in] HANDLE value);

    SetOutputArgumentOfArray(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfEnumeration(
        [in] Integer index,
        [in] Integer value);

    SetOutputArgumentOfEnumeration(
        [in] Integer index,
        [in] HANDLE addr);

    AssignOutputArgumentOfInterface(
        [in] Integer index,
        [in] IInterface* value);

    SetOutputArgumentOfInterface(
        [in] Integer index,
        [in] HANDLE addr);

    GetArgumentAddress(
        [in] Integer index,
        [out] HANDLE& addr);
}

}
