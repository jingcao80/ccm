//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {

[
    uuid(7eb63931-9e1d-4a39-b51f-a8e793aa98d7),
    version(0.1.0)
]
interface IMapEntry
{
    Equals(
        [in] IInterface* obj,
        [out] Boolean& result);

    GetHashCode(
        [out] Integer& hash);

    GetKey(
        [out] IInterface&& key);

    GetValue(
        [out] IInterface&& value);

    SetValue(
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);
}

interface ICollection;
interface ISet;

[
    uuid(76e49571-40d6-45f2-bb74-17045d67e64f),
    version(0.1.0)
]
interface IMap
{
    Clear();

    ContainsKey(
        [in] IInterface* key,
        [out] Boolean& result);

    ContainsValue(
        [in] IInterface* value,
        [out] Boolean& result);

    Equals(
        [in] IInterface* obj,
        [out] Boolean& result);

    Get(
        [in] IInterface* key,
        [out] IInterface&& value);

    GetEntrySet(
        [out] ISet&& entries);

    GetHashCode(
        [out] Integer& hash);

    GetKeySet(
        [out] ISet&& keys);

    GetSize(
        [out] Integer& size);

    GetValues(
        [out] ICollection&& values);

    IsEmpty(
        [out] Boolean& result);

    Put(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    PutAll(
        [in] IMap* m);

    PutIfAbsent(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    Remove(
        [in] IInterface* key,
        [out] IInterface** prevValue = nullptr);
}

}
}
