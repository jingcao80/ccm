//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::text::IDecimalFormatSymbols;
interface como::text::IFieldPosition;

namespace como {
namespace text {

/*
 * @Involve interface como::text::INumberFormat;
 * @Involve interface como::text::IFormat;
 * @Involve interface como::io::ISerializable;
 * @Involve interface como::core::ICloneable;
 */
[
    uuid(b1615f6c-db57-44fd-aa14-fd68dcc56992),
    version(0.1.0)
]
interface IDecimalFormat
{
    ApplyLocalizedPattern(
        [in] String pattern);

    ApplyPattern(
        [in] String pattern);

    GetDecimalFormatSymbols(
        [out] IDecimalFormatSymbols&& symbols);

    GetGroupingSize(
        [out] Integer& size);

    GetMultiplier(
        [out] Integer& multiplier);

    GetNegativePrefix(
        [out] String& prefix);

    GetNegativeSuffix(
        [out] String& suffix);

    GetPositivePrefix(
        [out] String& prefix);

    GetPositiveSuffix(
        [out] String& suffix);

    IsDecimalSeparatorAlwaysShown(
        [out] Boolean& shown);

    IsGroupingUsed(
        [out] Boolean& used);

    IsParseBigDecimal(
        [out] Boolean& value);

    IsParseIntegerOnly(
        [out] Boolean& value);

    SetDecimalFormatSymbols(
        [in] IDecimalFormatSymbols* symbols);

    SetDecimalSeparatorAlwaysShown(
        [in] Boolean shown);

    SetGroupingSize(
        [in] Integer size);

    SetGroupingUsed(
        [in] Boolean used);

    SetMultiplier(
        [in] Integer multiplier);

    SetNegativePrefix(
        [in] String prefix);

    SetNegativeSuffix(
        [in] String suffix);

    SetParseBigDecimal(
        [in] Boolean value);

    SetParseIntegerOnly(
        [in] Boolean value);

    SetPositivePrefix(
        [in] String prefix);

    SetPositiveSuffix(
        [in] String suffix);

    ToLocalizedPattern(
        [out] String& pattern);

    ToPattern(
        [out] String& pattern);
}

}
}
