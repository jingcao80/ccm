//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::util::IEnumeration;

namespace ccm {
namespace util {

/**
 * @Involve interface ccm::util::IList
 * @Involve interface ccm::util::ICollection
 * @Involve interface ccm::util::IRandomAccess
 * @Involve interface ccm::core::IIterable
 * @Involve interface ccm::core::ICloneable
 * @Involve interface ccm::io::ISerializable
 */
[
    uuid(496d3da5-9000-439e-bd01-3cf04a043f44),
    version(0.1.0)
]
interface IVector
{
    Add(
        [in] IInterface* e,
        [out] Boolean* changed = nullptr);

    Add(
        [in] Integer index,
        [in] IInterface* obj);

    AddAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    AddAll(
        [in] Integer index,
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    AddElement(
        [in] IInterface* e);

    Clear();

    Contains(
        [in] IInterface* obj,
        [out] Boolean* result);

    ContainsAll(
        [in] ICollection* c,
        [out] Boolean* result);

    CopyInto(
        [out] Array<IInterface*> anArray);

    EnsureCapacity(
        [in] Integer minCapacity);

    Get(
        [in] Integer index,
        [out] IInterface** obj);

    GetCapacity(
        [out] Integer* capacity);

    GetElementAt(
        [in] Integer index,
        [out] IInterface** element);

    GetElements(
        [out] IEnumeration** elements);

    GetFirstElement(
        [out] IInterface** element);

    GetIterator(
        [out] IIterator** it);

    GetLastElement(
        [out] IInterface** element);

    GetListIterator(
        [out] IListIterator** it);

    GetListIterator(
        [in] Integer index,
        [out] IListIterator** it);

    GetSize(
        [out] Integer* size);

    IndexOf(
        [in] IInterface* obj,
        [out] Integer* index);

    IndexOf(
        [in] IInterface* obj,
        [in] Integer fromIndex,
        [out] Integer* index);

    InsertElementAt(
        [in] IInterface* obj,
        [in] Integer index);

    IsEmpty(
        [out] Boolean* empty);

    LastIndexOf(
        [in] IInterface* obj,
        [out] Integer* index);

    LastIndexOf(
        [in] IInterface* obj,
        [in] Integer fromIndex,
        [out] Integer* index);

    Remove(
        [in] IInterface* obj,
        [out] Boolean* changed = nullptr);

    Remove(
        [in] Integer index,
        [out] IInterface** obj = nullptr);

    RemoveAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    RemoveAllElements();

    RemoveElement(
        [in] IInterface* obj,
        [out] Boolean* changed = nullptr);

    RemoveElementAt(
        [in] Integer index);

    RetainAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    Set(
        [in] Integer index,
        [in] IInterface* obj,
        [out] IInterface** prevObj = nullptr);

    SetElementAt(
        [in] IInterface* obj,
        [in] Integer index);

    SetSize(
        [in] Integer newSize);

    SubList(
        [in] Integer fromIndex,
        [in] Integer toIndex,
        [out] IList** subList);

    ToArray(
        [out, callee] Array<IInterface*>* objs);

    ToArray(
        [in] InterfaceID iid,
        [out, callee] Array<IInterface*>* objs);

    TrimToSize();
}

}
}
