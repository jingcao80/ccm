//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace io {

[
    uuid(6cac7adc-080b-417f-ab85-d0821bf88423),
    version(0.1.0)
]
interface IFloatBuffer
{
    AsReadOnlyBuffer(
        [out] IFloatBuffer** buffer);

    Compact();

    Duplicate(
        [out] IFloatBuffer** buffer);

    Get(
        [out] Float* f);

    Get(
        [in] Integer index,
        [out] Float* f);

    Get(
        [out] Array<Float>& dst);

    Get(
        [out] Array<Float>& dst,
        [in] Integer offset,
        [in] Integer length);

    GetOrder(
        [out] IByteOrder** bo);

    HasArray(
        [out] Boolean* result);

    Put(
        [in] Float f);

    Put(
        [in] Integer index,
        [in] Float f);

    Put(
        [in] Array<Float> src);

    Put(
        [in] Array<Float> src,
        [in] Integer offset,
        [in] Integer length);

    Put(
        [in] IFloatBuffer* src);

    Slice(
        [out] IFloatBuffer** buffer);
}

}
}
