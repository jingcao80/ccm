//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::util::ILocale;

namespace como {
namespace util {

[
    uuid(23187573-410c-46a8-b371-ebe00ab19fcc),
    version(0.1.0)
]
interface ICurrency
{
    GetCurrencyCode(
        [out] String* currency);

    GetDefaultFractionDigits(
        [out] Integer* digits);

    GetDisplayName(
        [out] String* displayName);

    GetDisplayName(
        [in] ILocale* locale,
        [out] String* displayName);

    GetNumericCode(
        [out] Integer* numericCode);

    GetSymbol(
        [out] String* symbol);

    GetSymbol(
        [in] ILocale* locale,
        [out] String* symbol);
}

}
}
