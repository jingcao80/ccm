//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::util::IMapEntry;

namespace como {
namespace util {

/**
 * @Involve interface como::util::IMap
 * @Involve interface como::core::ICloneable
 * @Involve interface como::io::ISerializable
 */
[
    uuid(b916c8bb-1d3e-4c7b-9d68-794c586a5e46),
    version(0.1.0)
]
interface ILinkedHashMap
{
    GetEldest(
        [out] IMapEntry&& entry);
}

}
}
