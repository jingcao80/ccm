//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {
namespace concurrent {

/*
 * @Involve interface ccm::util::IRandom
 */
[
    uuid(100a074a-b631-4d9f-80a8-f83c67655f5a),
    version(0.1.0)
]
interface IThreadLocalRandom
{
    NextDouble(
        [in] Double bound,
        [out] Double* value);

    NextDouble(
        [in] Double origin,
        [in] Double bound,
        [out] Double* value);

    NextInt(
        [in] Integer origin,
        [in] Integer bound,
        [out] Integer* value);

    NextLong(
        [in] Long bound,
        [out] Long* value);

    NextLong(
        [in] Long origin,
        [in] Long bound,
        [out] Long* value);
}

}
}
}
