//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace io {

/*
 * @involve como::io::ICloseable
 * @involve como::core::IAutoCloseable
 * @involve como::io::IFlushable
 */
[
    uuid(46274ade-a4d4-4200-8d95-59b40160cf68),
    version(0.1.0)
]
interface IOutputStream
{
    Close();

    Flush();

    Write(
        [in] Integer byte);

    Write(
        [in] Array<Byte> buffer);

    Write(
        [in] Array<Byte> buffer,
        [in] Integer offset,
        [in] Integer size);
}

}
}
