//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {

interface IMetaMethod;
interface IArgumentList;

[
    uuid(bf89f2ce-ba5f-4f5d-a866-9e34048ee009),
    version(0.1.0)
]
interface IInvocationHandler
{
    Invoke(
        [in] IInterface* proxy,
        [in] IMetaMethod* method,
        [in] IArgumentList* args);
}

interface IDeathRecipient;

[
    uuid(2598f97d-0e6b-45a2-8c21-ffeca8347233),
    version(0.1.0)
]
interface IProxy
{
    SetInvocationHandler(
        [in] IInvocationHandler* handler);

    IsStubAlive(
        [out] Boolean* alive);

    LinkToDeath(
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0);

    UnlinkToDeath(
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0,
        [out] IDeathRecipient** outRecipient = nullptr);
}

[
    uuid(2598f97d-0e6b-45a2-8c21-ffeca8347233),
    version(0.1.0)
]
interface IDeathRecipient
{
    ProxyDied(
        [out] IProxy** who);
}

[
    uuid(7752e566-880a-4abd-99b9-417176e0644f),
    version(0.1.0)
]
interface IStub
{
    Invoke(
        [in] IMetaMethod* method,
        [in] IArgumentList* args);
}

}
