//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::security::IProvider;

namespace ccm {
namespace security {
namespace cca {

[
    uuid(2c685889-e192-41fe-953b-2dbffc54203a),
    version(0.1.0)
]
interface IInstance
{
    GetImpl(
        [out] IInterface** impl);

    GetProvider(
        [out] IProvider** provider);
}

[
    uuid(b8e28501-8a94-4767-b5e9-60e6793f49f8),
    version(0.1.0)
]
interface IInstanceFactory
{}

}
}
}
