//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {

/**
 * @Involve interface ccm::util::IList
 * @Involve interface ccm::util::ICollection
 * @Involve interface ccm::util::IRandomAccess
 * @Involve interface ccm::core::IIterable
 * @Involve interface ccm::core::ICloneable
 * @Involve interface ccm::io::ISerializable
 */
[
    uuid(496d3da5-9000-439e-bd01-3cf04a043f44),
    version(0.1.0)
]
interface IVector
{
    Add(
        [in] IInterface* e,
        [out] Boolean* changed = nullptr);

    AddElement(
        [in] IInterface* e);

    ElementAt(
        [in] Integer index,
        [out] IInterface** obj);

    Get(
        [in] Integer index,
        [out] IInterface** obj);

    GetSize(
        [out] Integer* size);

    IndexOf(
        [in] IInterface* obj,
        [out] Integer* index);

    Set(
        [in] Integer index,
        [in] IInterface* obj,
        [out] IInterface** prevObj = nullptr);

    SetSize(
        [in] Integer newSize);
}

}
}
