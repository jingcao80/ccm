//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ccm/core/Errors.cdl"
include "ccm/core/Exceptions.cdl"
include "ccm/core/IAnnotation.cdl"
include "ccm/core/IAppendable.cdl"
include "ccm/core/IArray.cdl"
include "ccm/core/IArrayHolder.cdl"
include "ccm/core/IAutoCloseable.cdl"
include "ccm/core/IBoolean.cdl"
include "ccm/core/IByte.cdl"
include "ccm/core/IChar.cdl"
include "ccm/core/ICharSequence.cdl"
include "ccm/core/ICloneable.cdl"
include "ccm/core/IComparable.cdl"
include "ccm/core/IDouble.cdl"
include "ccm/core/IFloat.cdl"
include "ccm/core/IInteger.cdl"
include "ccm/core/IIterable.cdl"
include "ccm/core/ILong.cdl"
include "ccm/core/INumber.cdl"
include "ccm/core/IReadable.cdl"
include "ccm/core/IRunnable.cdl"
include "ccm/core/IRuntime.cdl"
include "ccm/core/ISecurityManager.cdl"
include "ccm/core/IShort.cdl"
include "ccm/core/IStackTrace.cdl"
include "ccm/core/IStackTraceElement.cdl"
include "ccm/core/IString.cdl"
include "ccm/core/IStringBuffer.cdl"
include "ccm/core/IStringBuilder.cdl"
include "ccm/core/ISynchronize.cdl"
include "ccm/core/ISystem.cdl"
include "ccm/core/IThread.cdl"
include "ccm/core/IThreadGroup.cdl"
include "ccm/core/IThreadLocal.cdl"

namespace ccm {
namespace core {

[
    uuid(bc5be123-34ab-4373-ab98-31c3e3c68b1b),
    version(0.1.0)
]
coclass CArray
{
    Constructor(
        [in] InterfaceID elemId,
        [in] Long size);

    interface IArray;
}

[
    uuid(f608b0cd-d0af-4adb-a2a4-6f241136b992),
    version(0.1.0)
]
coclass CArrayHolder
{
    Constructor(
        [in] Triple array);

    interface IArrayHolder;
}

[
    uuid(6cdec0e6-ee66-4ba3-b167-e8d45e029fbd),
    version(0.1.0)
]
coclass CSystem
{
    interface ISystem;
}

[
    uuid(339a8069-7448-4d12-9c50-d45497fb245b),
    version(0.1.0)
]
coclass CThread
{
    Constructor();

    Constructor(
        [in] IThreadGroup* group,
        [in] String name,
        [in] Integer priority,
        [in] Boolean daemon);

    // @hide
    Constructor(
        [in] HANDLE peer);

    interface IRunnable;
    interface IThread;
}

[
    uuid(730c7375-05c3-4b86-933c-ab2808164280),
    version(0.1.0)
]
coclass CThreadGroup
{
    // @hide
    Constructor();

    Constructor(
        [in] String name);

    Constructor(
        [in] IThreadGroup* parent,
        [in] String name);

    interface IThreadGroup;
}

[
    uuid(dce1a0c3-b23d-4b89-bdaf-8a1bf581ee44),
    version(0.1.0)
]
coclass CThreadLocal
{
    Constructor();

    interface IThreadLocal;
}

}
}
