//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace io {

[
    uuid(73dcfab7-ea7a-4bab-af32-4c3d0ad6b986),
    version(0.1.0)
]
interface IBuffer
{
    Clear();

    Flip();

    GetArray(
        [out, callee] Array<IInterface*>* array);

    GetArrayOffset(
        [out] Integer* offset);

    GetCapacity(
        [out] Integer* capacity);

    GetLimit(
        [out] Integer* limit);

    GetPosition(
        [out] Integer* position);

    HasArray(
        [out] Boolean* result);

    HasRemaining(
        [out] Boolean* result);

    IsDirect(
        [out] Boolean* direct);

    IsReadOnly(
        [out] Boolean* readOnly);

    Mark();

    Remaining(
        [out] Integer* remaining);

    Reset();

    Rewind();

    SetLimit(
        [in] Integer newLimit);

    SetPosition(
        [in] Integer newPosition);
}

}
}
