//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {
namespace concurrent {

/*
 * @Involve interface como::util::IRandom
 * @Involve interface como::io:ISerializable
 */
[
    uuid(100a074a-b631-4d9f-80a8-f83c67655f5a),
    version(0.1.0)
]
interface IThreadLocalRandom
{
    NextDouble(
        [in] Double bound,
        [out] Double* value);

    NextDouble(
        [in] Double origin,
        [in] Double bound,
        [out] Double* value);

    NextInteger(
        [in] Integer origin,
        [in] Integer bound,
        [out] Integer* value);

    NextLong(
        [in] Long bound,
        [out] Long* value);

    NextLong(
        [in] Long origin,
        [in] Long bound,
        [out] Long* value);
}

}
}
}
