//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace security {

/*
 * @Involve interface ccm::util::IProperties;
 * @Involve interface ccm::util::IHashtable;
 * @Involve interface ccm::util::IDictionary;
 * @Involve interface ccm::util::IMap;
 * @Involve interface ccm::core::ICloneable;
 * @Involve interface ccm::io::ISerializable;
 */
[
    uuid(5175ea7f-5a2b-480e-b8c5-37bef4036c6a),
    version(0.1.0)
]
interface IProvider
{}

}
}
