//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::core::IStringBuffer;
interface como::text::IAttributedCharacterIterator;
interface como::text::IFieldPosition;
interface como::text::IParsePosition;
interface como::util::ILocale;

namespace como {
namespace text {

/**
 * @Involve interface como::text::IFormatField
 */
[
    uuid(484a7e85-38ac-427a-b6b6-2ec6e6d51176),
    version(0.1.0)
]
interface IMessageFormatField {
}

/*
 * @Involve interface como::text::IFormat;
 * @Involve interface como::io::ISerializable;
 * @Involve interface como::core::ICloneable;
 */
[
    uuid(207d608f-1ca5-4ae1-8723-b36e26f25048),
    version(0.1.0)
]
interface IMessageFormat
{
    ApplyPattern(
        [in] String pattern);

    Format(
        [in] Array<IInterface*> arguments,
        [out] IStringBuffer* result,
        [in] IFieldPosition* pos);

    Format(
        [in] IInterface* arguments,
        [in] IStringBuffer* result,
        [in] IFieldPosition* pos);

    FormatToCharacterIterator(
        [in] IInterface* arguments,
        [out] IAttributedCharacterIterator** cit);

    GetFormats(
        [out, callee] Array<IFormat*>* formats);

    GetFormatsByArgumentIndex(
        [out, callee] Array<IFormat*>* formats);

    GetLocale(
        [out] ILocale** locale);

    Parse(
        [in] String source,
        [out, callee] Array<IInterface*>* result);

    Parse(
        [in] String source,
        [in] IParsePosition* pos,
        [out, callee] Array<IInterface*>* result);

    ParseObject(
        [in] String source,
        [in] IParsePosition* pos,
        [out] IInterface** result);

    SetFormat(
        [in] Integer formatElementIndex,
        [in] IFormat* newFormat);

    SetFormatByArgumentIndex(
        [in] Integer argumentIndex,
        [in] IFormat* newFormat);

    SetFormats(
        [in] Array<IFormat*> newFormats);

    SetFormatsByArgumentIndex(
        [in] Array<IFormat*> newFormats);

    SetLocale(
        [in] ILocale* locale);

    ToPattern(
        [out] String* pattern);
}

}
}
