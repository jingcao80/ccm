//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {

enum RPCType
{
    Local,
    Remote
}

enum RPCPeer
{
    Proxy,
    Stub
}

[
    uuid(3d29cb55-f7d1-4b79-9e63-ad14a57fd9f1),
    version(0.1.0)
]
interface IParcel
{
    ReadChar(
        [out] Char* value);

    WriteChar(
        [in] Char value);

    ReadByte(
        [out] Byte* value);

    WriteByte(
        [in] Byte value);

    ReadShort(
        [out] Short* value);

    WriteShort(
        [in] Short value);

    ReadInteger(
        [out] Integer* value);

    WriteInteger(
        [in] Integer value);

    ReadLong(
        [out] Long* value);

    WriteLong(
        [in] Long value);

    ReadFloat(
        [out] Float* value);

    WriteFloat(
        [in] Float value);

    ReadDouble(
        [out] Double* value);

    WriteDouble(
        [in] Double value);

    ReadBoolean(
        [out] Boolean* value);

    WriteBoolean(
        [in] Boolean value);

    ReadString(
        [out] String* value);

    WriteString(
        [in] String value);

    ReadCoclassID(
        [out] CoclassID* value);

    WriteCoclassID(
        [in] CoclassID value);

    ReadComponentID(
        [out] ComponentID* value);

    WriteComponentID(
        [in] ComponentID value);

    ReadInterfaceID(
        [out] InterfaceID* value);

    WriteInterfaceID(
        [in] InterfaceID value);

    ReadECode(
        [out] ECode* value);

    WriteECode(
        [in] ECode value);

    ReadEnumeration(
        [out] Integer* value);

    WriteEnumeration(
        [in] Integer value);

    ReadArray(
        [out] HANDLE array);

    WriteArray(
        [in] HANDLE array);

    ReadInterface(
        [out] IInterface** value);

    WriteInterface(
        [in] IInterface* value);

    GetDataPayload(
        [out] HANDLE* data);

    GetDataSize(
        [out] Long* size);

    SetDataPosition(
        [in] Long pos);
}

interface IArgumentList;
interface IDeathRecipient;
interface IMetaMethod;
interface IProxy;

[
    uuid(bf89f2ce-ba5f-4f5d-a866-9e34048ee009),
    version(0.1.0)
]
interface IRPCChannel
{
    GetRPCType(
        [out] RPCType* type);

    CreateArgumentParcel(
        [out] IParcel** parcel);

    IsPeerAlive(
        [out] Boolean* alive);

    LinkToDeath(
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0);

    UnlinkToDeath(
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0,
        [out] IDeathRecipient** outRecipient = nullptr);

    Invoke(
        [in] IProxy* proxy,
        [in] IMetaMethod* method,
        [in] IParcel* argParcel,
        [out] IParcel** resParcel);

    StartListening();
}

[
    uuid(d1adf1f9-2062-45fd-aa33-edd481a04417),
    version(0.1.0)
]
interface IRPCChannelFactory
{
    CreateChannel(
        [in] RPCPeer peer,
        [out] IRPCChannel** channel);
}

[
    uuid(2598f97d-0e6b-45a2-8c21-ffeca8347233),
    version(0.1.0)
]
interface IProxy
{
    GetTargetCoclass(
        [out] IMetaCoclass** target);

    IsStubAlive(
        [out] Boolean* alive);

    LinkToDeath(
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0);

    UnlinkToDeath(
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0,
        [out] IDeathRecipient** outRecipient = nullptr);
}

[
    uuid(2598f97d-0e6b-45a2-8c21-ffeca8347233),
    version(0.1.0)
]
interface IDeathRecipient
{
    ProxyDied(
        [out] IProxy** who);
}

[
    uuid(7752e566-880a-4abd-99b9-417176e0644f),
    version(0.1.0)
]
interface IStub
{
    Invoke(
        [in] IMetaMethod* method,
        [in] IArgumentList* args);
}

}
