//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::IMetaCoclass;
interface ccm::IMetaComponent;

namespace ccm {

[
    uuid(00000000-0000-0000-0000-000000000002),
    version(0.1.0)
]
interface IClassObject
{
    AttachMetadata(
        [in] IMetaComponent* component);

    CreateObject(
        [in] InterfaceID iid,
        [out] IInterface** object);
}

[
    uuid(00000000-0000-0000-0000-000000000003),
    version(0.1.0)
]
interface IObject
{
    AttachMetadata(
        [in] IMetaComponent* component,
        [in] String coclassName);

    GetCoclassID(
        [out] CoclassID* cid);

    GetCoclass(
        [out] IMetaCoclass** klass);

    GetHashCode(
        [out] Integer* hash);

    Equals(
        [in] IInterface* obj,
        [out] Boolean* same);

    ToString(
        [out] String* desc);
}

[
    uuid(00000000-0000-0000-0000-000000000004),
    version(0.1.0)
]
interface IClassLoader
{
    LoadComponent(
        [in] ComponentID compId,
        [out] IMetaComponent** component);

    UnloadComponent(
        [in] ComponentID compId);

    LoadCoclass(
        [in] String fullName,
        [out] IMetaCoclass** klass);
}

[
    uuid(00000000-0000-0000-0000-000000000005),
    version(0.1.0)
]
interface IWeakReference
{
    Resolve(
        [in] InterfaceID iid,
        [out] IInterface** object);
}

[
    uuid(00000000-0000-0000-0000-000000000006),
    version(0.1.0)
]
interface IWeakReferenceSource
{
    GetWeakReference(
        [out] IWeakReference** wr);
}

}
