//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ccm/misc/IFDBigInteger.cdl"
include "ccm/misc/IFloatingDecimal.cdl"
include "ccm/misc/IFormattedFloatingDecimal.cdl"

namespace ccm {
namespace misc {

[
    uuid(e8cd20cc-761f-4006-9741-fe8cf701c009),
    version(0.1.0)
]
coclass CFDBigInteger
{
    Constructor(
        [in] Long lValue,
        [in] Array<Char> digits,
        [in] Integer kDigits,
        [in] Integer nDigits);

    interface IFDBigInteger;
}

}
}
