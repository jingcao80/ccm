//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "como/io/Errors.cdl"
include "como/io/Exceptions.cdl"
include "como/io/IBuffer.cdl"
include "como/io/IBufferedWriter.cdl"
include "como/io/IByteArrayOutputStream.cdl"
include "como/io/IByteBuffer.cdl"
include "como/io/IByteOrder.cdl"
include "como/io/ICharBuffer.cdl"
include "como/io/ICloseable.cdl"
include "como/io/IDataInput.cdl"
include "como/io/IDoubleBuffer.cdl"
include "como/io/IFile.cdl"
include "como/io/IFileDescriptor.cdl"
include "como/io/IFileFilter.cdl"
include "como/io/IFileInputStream.cdl"
include "como/io/IFileOutputStream.cdl"
include "como/io/IFilenameFilter.cdl"
include "como/io/IFloatBuffer.cdl"
include "como/io/IFlushable.cdl"
include "como/io/IInputStream.cdl"
include "como/io/IIntegerBuffer.cdl"
include "como/io/IInterruptible.cdl"
include "como/io/ILongBuffer.cdl"
include "como/io/IMappedByteBuffer.cdl"
include "como/io/IObjectInput.cdl"
include "como/io/IObjectInputStream.cdl"
include "como/io/IOutputStream.cdl"
include "como/io/IOutputStreamWriter.cdl"
include "como/io/IPrintStream.cdl"
include "como/io/IPrintWriter.cdl"
include "como/io/IReader.cdl"
include "como/io/ISerializable.cdl"
include "como/io/IShortBuffer.cdl"
include "como/io/IStringWriter.cdl"
include "como/io/IWriter.cdl"
include "como/io/channels/IDirectBuffer.cdl"
include "como/io/channels/IFileChannel.cdl"
include "como/io/charset/ICharset.cdl"
include "como/io/charset/ICharsetDecoder.cdl"
include "como/io/charset/ICharsetEncoder.cdl"
include "como/io/charset/ICodingErrorAction.cdl"
include "como/io/charset/ICoderResult.cdl"
include "como/io/charset/IStreamEncoder.cdl"
include "como/io/charset/spi/ICharsetProvider.cdl"

interface como::core::IAppendable;
interface como::core::IAutoCloseable;
interface como::core::IComparable;
interface como::io::channels::IDirectBuffer;
interface como::io::charset::ICharset;
interface como::io::charset::ICharsetEncoder;
interface como::net::IURI;

namespace como {
namespace io {

[
    uuid(cf7b3ffb-46ce-44fc-9057-d8ec03c820b7),
    version(0.1.0)
]
coclass CBufferedWriter
{
    Constructor(
        [in] IWriter* outW);

    Constructor(
        [in] IWriter* outW,
        [in] Integer sz);

    interface IBufferedWriter;
    interface IWriter;
    interface IAppendable;
    interface ICloseable;
    interface IFlushable;
    interface IAutoCloseable;
}

[
    uuid(69455e4d-56b1-43b1-98b1-e4907e332a4f),
    version(0.1.0)
]
coclass CByteArrayOutputStream
{
    Constructor();

    Constructor(
        [in] Integer size);

    interface IByteArrayOutputStream;
    interface IOutputStream;
    interface IFlushable;
    interface ICloseable;
    interface IAutoCloseable;
}

[
    uuid(160997fd-1165-46dd-a47a-8a000bcd1916),
    version(0.1.0)
]
coclass CDirectByteBuffer
{
    Constructor(
        [in] Integer cap,
        [in] HANDLE address,
        [in] IFileDescriptor* fd,
        [in] Boolean isReadOnly);

    interface IDirectBuffer;
    interface IMappedByteBuffer;
    interface IByteBuffer;
    interface IBuffer;
    interface IComparable;
}

[
    uuid(0d9c5571-7eaa-44e1-815f-c6af421c780d),
    version(0.1.0)
]
coclass CFile
{
    Constructor(
        [in] String pathname);

    Constructor(
        [in] String parent,
        [in] String child);

    Constructor(
        [in] IFile* parent,
        [in] String child);

    Constructor(
        [in] IURI* urii);

    // @hide
    Constructor(
        [in] String pathname,
        [in] Integer prefixLength);

    // @hide
    Constructor(
        [in] String child,
        [in] IFile* parent);

    interface IFile;
}

[
    uuid(3e291dd3-0c31-4526-8ef9-fe61bc1e508e),
    version(0.1.0)
]
coclass CFileDescriptor
{
    Constructor();

    Constructor(
        [in] Integer descriptor);

    interface IFileDescriptor;
}

[
    uuid(28063bc3-48b2-43f4-b159-c4c65475b844),
    version(0.1.0)
]
coclass CFileInputStream
{
    Constructor(
        [in] String name);

    Constructor(
        [in] IFile* file);

    Constructor(
        [in] IFileDescriptor* fdObj);

    Constructor(
        [in] IFileDescriptor* fdObj,
        [in] Boolean isFdOwner);

    interface IFileInputStream;
    interface IInputStream;
    interface ICloseable;
    interface IAutoCloseable;
}

[
    uuid(6d5f9b98-ce5c-4e30-a5ca-c0c74e0dc8fd),
    version(0.1.0)
]
coclass CFileOutputStream
{
    Constructor(
        [in] String name);

    Constructor(
        [in] String name,
        [in] Boolean append);

    Constructor(
        [in] IFile* file);

    Constructor(
        [in] IFile* file,
        [in] Boolean append);

    Constructor(
        [in] IFileDescriptor* fdObj);

    Constructor(
        [in] IFileDescriptor* fdObj,
        [in] Boolean isFdOwner);

    interface IFileOutputStream;
    interface IOutputStream;
    interface IFlushable;
    interface ICloseable;
    interface IAutoCloseable;
}

[
    uuid(3f1442a5-ce76-40b3-8889-c9431c810c1d),
    version(0.1.0)
]
coclass COutputStreamWriter
{
    Constructor(
        [in] IOutputStream* outstream,
        [in] String charsetName);

    Constructor(
        [in] IOutputStream* outstream);

    Constructor(
        [in] IOutputStream* outstream,
        [in] ICharset* cs);

    Constructor(
        [in] IOutputStream* outstream,
        [in] ICharsetEncoder* enc);

    interface IOutputStreamWriter;
    interface IWriter;
    interface IAppendable;
    interface ICloseable;
    interface IFlushable;
    interface IAutoCloseable;
}

[
    uuid(5de87670-f240-43cd-b06d-a758b4914e76),
    version(0.1.0)
]
coclass CPrintWriter
{
    Constructor(
        [in] IWriter* outstream);

    Constructor(
        [in] IWriter* outstream,
        [in] Boolean autoFlush);

    Constructor(
        [in] IOutputStream* outstream);

    Constructor(
        [in] IOutputStream* outstream,
        [in] Boolean autoFlush);

    Constructor(
        [in] String fileName);

    Constructor(
        [in] String fileName,
        [in] String csn);

    Constructor(
        [in] IFile* file);

    Constructor(
        [in] IFile* file,
        [in] String csn);

    interface IPrintWriter;
}

[
    uuid(2a886435-1ec8-4311-be20-03cff45b0dc8),
    version(0.1.0)
]
coclass CStringWriter
{
    Constructor();

    Constructor(
        [in] Integer initialSize);

    interface IStringWriter;
    interface IWriter;
    interface IAppendable;
    interface ICloseable;
    interface IFlushable;
    interface IAutoCloseable;
}

}
}
