//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::math::IBigDecimal;

namespace ccm {
namespace math {

enum RoundingMode {
    /**
     * Rounding mode where positive values are rounded towards positive infinity
     * and negative values towards negative infinity.
     * Rule: {x.round().abs() >= x.abs()}
     */
    UP = IBigDecimal::ROUND_UP,

    /**
     * Rounding mode where the values are rounded towards zero.
     * Rule: {x.round().abs() <= x.abs()}
     */
    DOWN = IBigDecimal::ROUND_DOWN,

    /**
     * Rounding mode to round towards positive infinity. For positive values
     * this rounding mode behaves as {#UP}, for negative values as
     * {#DOWN}.
     * Rule: {x.round() >= x}
     */
    CEILING = IBigDecimal::ROUND_CEILING,

    /**
     * Rounding mode to round towards negative infinity. For positive values
     * this rounding mode behaves as {#DOWN}, for negative values as
     * {#UP}.
     * Rule: {x.round() <= x}
     */
    FLOOR = IBigDecimal::ROUND_FLOOR,

    /**
     * Rounding mode where values are rounded towards the nearest neighbor. Ties
     * are broken by rounding up.
     */
    HALF_UP = IBigDecimal::ROUND_HALF_UP,

    /**
     * Rounding mode where values are rounded towards the nearest neighbor. Ties
     * are broken by rounding down.
     */
    HALF_DOWN = IBigDecimal::ROUND_HALF_DOWN,

    /**
     * Rounding mode where values are rounded towards the nearest neighbor. Ties
     * are broken by rounding to the even neighbor.
     */
    HALF_EVEN = IBigDecimal::ROUND_HALF_EVEN,

    /**
     * Rounding mode where the rounding operations throws an ArithmeticException
     * for the case that rounding is necessary, i.e. for the case that the value
     * cannot be represented exactly.
     */
    UNNECESSARY = IBigDecimal::ROUND_UNNECESSARY
}

}
}
