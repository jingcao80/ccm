//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {

interface IEnumeration;

[
    uuid(6e0f6eb5-6c0e-4f31-b042-d5cd18cf8a23),
    version(0.1.0)
]
interface IDictionary
{
    Get(
        [in] IInterface* key,
        [out] IInterface&& value);

    GetElements(
        [out] IEnumeration&& elements);

    GetKeys(
        [out] IEnumeration&& keys);

    GetSize(
        [out] Integer& size);

    IsEmpty(
        [out] Boolean& result);

    Put(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    Remove(
        [in] IInterface* key,
        [out] IInterface** prevValue = nullptr);
}

}
}
