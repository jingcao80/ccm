//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace core {

[
    uuid(9549d2b9-6356-42fa-92bd-5d8ea657e5e6),
    version(0.1.0)
]
interface IArrayHolder
{
    const Integer TYPE_UNKNOWN_ARRAY = 0;

    const Integer TYPE_CHAR_ARRAY = 1;

    const Integer TYPE_BYTE_ARRAY = 2;

    const Integer TYPE_SHORT_ARRAY = 3;

    const Integer TYPE_INTEGER_ARRAY = 4;

    const Integer TYPE_LONG_ARRAY = 5;

    const Integer TYPE_FLOAT_ARRAY = 6;

    const Integer TYPE_DOUBLE_ARRAY = 7;

    const Integer TYPE_BOOLEAN_ARRAY = 8;

    const Integer TYPE_STRING_ARRAY = 9;

    const Integer TYPE_INTERFACE_ARRAY = 17;

    GetArray(
        [out] Triple* array);

    GetArrayType(
        [out] Integer& type);
}

}
}
