//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::core::IInteger;
interface como::core::ILong;
interface como::util::ITimeZone;
interface como::util::calendar::IEra;

namespace como {
namespace util {
namespace calendar {

/*
 * @Involve interface como::core::ICloneable
 */
[
    uuid(251aa366-dca8-48c5-b0d7-27a33657ae75),
    version(0.1.0)
]
interface ICalendarDate
{
    const Integer FIELD_UNDEFINED = IInteger::MIN_VALUE;

    const Long TIME_UNDEFINED = ILong::MIN_VALUE;

    AddDate(
        [in] Integer year,
        [in] Integer month,
        [in] Integer dayOfMonth);

    AddDayOfMonth(
        [in] Integer n);

    AddHours(
        [in] Integer n);

    AddMillis(
        [in] Integer n);

    AddMinutes(
        [in] Integer n);

    AddMonth(
        [in] Integer n);

    AddSeconds(
        [in] Integer n);

    AddTimeOfDay(
        [in] Integer hours,
        [in] Integer minutes,
        [in] Integer seconds,
        [in] Integer millis);

    AddYear(
        [in] Integer n);

    GetDaylightSaving(
        [out] Integer* ds);

    GetDayOfMonth(
        [out] Integer* date);

    GetDayOfWeek(
        [out] Integer* date);

    GetEra(
        [out] IEra** era);

    GetHours(
        [out] Integer* hours);

    GetMillis(
        [out] Integer* millis);

    GetMinutes(
        [out] Integer* minutes);

    GetMonth(
        [out] Integer* month);

    GetSeconds(
        [out] Integer* seconds);

    GetTimeOfDay(
        [out] Long* date);

    GetYear(
        [out] Integer* year);

    GetZone(
        [out] ITimeZone** zone);

    GetZoneOffset(
        [out] Integer* offset);

    IsDaylightTime(
        [out] Boolean* daylightTime);

    IsLeapYear(
        [out] Boolean* leapYear);

    IsNormalized(
        [out] Boolean* normalized);

    IsSameDate(
        [in] ICalendarDate* date,
        [out] Boolean* same);

    IsStandardTime(
        [out] Boolean* standardTime);

    SetDate(
        [in] Integer year,
        [in] Integer month,
        [in] Integer dayOfMonth);

    SetDaylightSaving(
        [in] Integer daylightSaving);

    SetDayOfMonth(
        [in] Integer date);

    SetDayOfWeek(
        [in] Integer dayOfWeek);

    SetEra(
        [in] IEra* era);

    SetHours(
        [in] Integer hours);

    SetLeapYear(
        [in] Boolean leapYear);

    SetMillis(
        [in] Integer millis);

    SetMinutes(
        [in] Integer minutes);

    SetMonth(
        [in] Integer month);

    SetNormalized(
        [in] Boolean normalized);

    SetSeconds(
        [in] Integer seconds);

    SetStandardTime(
        [in] Boolean standardTime);

    SetTimeOfDay(
        [in] Long fraction);

    SetTimeOfDay(
        [in] Integer hours,
        [in] Integer minutes,
        [in] Integer seconds,
        [in] Integer millis);

    SetYear(
        [in] Integer year);

    SetZone(
        [in] ITimeZone* zoneinfo);

    SetZoneOffset(
        [in] Integer offset);
}

}
}
}
