//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

[
    uuid(6a07eff9-9090-41a9-bfc3-67eb3ed80f49),
    url("http://ccm.org/component/sample/FooBarDemo.so")
]
module FooBarDemo
{

include "IFoo.cdl"
include "IBar.cdl"

namespace ccm {
namespace demo {

[
    uuid(b150ddc0-530b-411f-8462-b04252fd012b),
    version(0.1.0)
]
coclass CFoo
{
    interface IFoo;
}

[
    uuid(855db520-7f7a-4ad1-a60a-7d8d3461be7b),
    version(0.1.0)
]
coclass CFooBar
{
    constructor();

    constructor(
        [in] Long data);

    interface IFoo;
    interface IBar;
}

}
}

}
