//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {

interface IMap;
interface ISet;

[
    uuid(b60ce103-12d2-4b1f-ae56-b5d5feec23d2),
    version(0.1.0)
]
interface IHashtable
{
    Clear();

    Contains(
        [in] IInterface* value,
        [out] Boolean& result);

    ContainsKey(
        [in] IInterface* key,
        [out] Boolean& result);

    ContainsValue(
        [in] IInterface* value,
        [out] Boolean& result);

    Equals(
        [in] IInterface* obj,
        [out] Boolean& result);

    Get(
        [in] IInterface* key,
        [out] IInterface&& value);

    GetElements(
        [out] IEnumeration&& elements);

    GetEntrySet(
        [out] ISet&& entries);

    GetHashCode(
        [out] Integer& hash);

    GetKeys(
        [out] IEnumeration&& keys);

    GetValues(
        [out] ICollection&& values);

    GetKeySet(
        [out] ISet&& keys);

    GetSize(
        [out] Integer& size);

    IsEmpty(
        [out] Boolean& result);

    Put(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    PutAll(
        [in] IMap* m);

    Remove(
        [in] IInterface* key,
        [out] IInterface** prevValue = nullptr);
}

}
}
