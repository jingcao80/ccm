//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::io::IFile;

namespace como {
namespace io {

[
    uuid(5135c5a7-1174-430b-93f6-548b17a436cf),
    version(0.1.0)
]
interface IFileFilter
{
    Accept(
        [in] IFile* pathname,
        [out] Boolean& accepted);
}

}
}
