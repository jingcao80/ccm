//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::util::IIterator;

namespace ccm {
namespace util {

/*
 * @Involve interface ccm::util::ISet
 * @Involve interface ccm::util::ICollection
 * @Involve interface ccm::io::ISerializable
 * @Involve interface ccm::core::IIterable
 * @Involve interface ccm::core::ICloneable
 */
[
    uuid(4f2e0d90-13b0-4ac9-857a-caaf328e4216),
    version(0.1.0)
]
interface IHashSet
{
    Add(
        [in] IInterface* obj,
        [out] Boolean* modified = nullptr);

    AddAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    Clear();

    Contains(
        [in] IInterface* obj,
        [out] Boolean* result);

    ContainsAll(
        [in] ICollection* c,
        [out] Boolean* result);

    Equals(
        [in] IInterface* obj,
        [out] Boolean* result);

    GetHashCode(
        [out] Integer* hash);

    GetIterator(
        [out] IIterator** it);

    GetSize(
        [out] Integer* size);

    IsEmpty(
        [out] Boolean* result);

    Remove(
        [in] IInterface* obj,
        [out] Boolean* contained = nullptr);

    RemoveAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    RetainAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    ToArray(
        [out, callee] Array<IInterface*>* objs);

    ToArray(
        [in] InterfaceID iid,
        [out, callee] Array<IInterface*>* objs);
}

}
}
