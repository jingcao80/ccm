//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace text {

/*
 * @Involve interface ccm::io::ISerializable
 * @Involve interface ccm::core::ICloneable
 */
[
    uuid(b2e89609-5020-4f1a-ae3b-3406c4021da1),
    version(0.1.0)
]
interface IDateFormatSymbols
{
    GetAmPmStrings(
        [out, callee] Array<String>* ampm);

    GetEras(
        [out, callee] Array<String>* eras);

    GetMonths(
        [out, callee] Array<String>* months);

    GetShortMonths(
        [out, callee] Array<String>* months);

    GetShortWeekdays(
        [out, callee] Array<String>* weekdays);

    GetWeekdays(
        [out, callee] Array<String>* weekdays);
}

}
}
