//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace io {

const Integer E_IO_EXCEPTION = 0x80010300;
const Integer E_IO_SYNC_FAILED_EXCEPTION = 0x80010301;
const Integer E_FILE_NOT_FOUND_EXCEPTION = 0x80010302;
const Integer E_USE_MANUAL_SKIP_EXCEPTION = 0x80010303;
const Integer E_INTERRUPTED_IO_EXCEPTION = 0x80010304;
const Integer E_UNSUPPORTED_ENCODING_EXCEPTION = 0x80010305;
const Integer E_INVALID_OBJECT_EXCEPTION = 0x80010306;
const Integer E_INVALID_MARK_EXCEPTION = 0x80010307;
const Integer E_BUFFER_UNDERFLOW_EXCEPTION = 0x80010308;
const Integer E_BUFFER_OVERFLOW_EXCEPTION = 0x80010309;
const Integer E_READ_ONLY_BUFFER_EXCEPTION = 0x8001030a;
const Integer E_UNSUPPORTED_CHARSET_EXCEPTION = 0x8001030b;
const Integer E_ILLEGAL_CHARSET_NAME_EXCEPTION = 0x8001030c;
const Integer E_MALFORMED_INPUT_EXCEPTION = 0x8001030d;
const Integer E_UNMAPPABLE_CHARACTER_EXCEPTION = 0x8001030e;

}
}
