//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace io {

/*
 * @Involve interface ccm::io::IBuffer;
 * @Involve interface ccm::core::IComparable;
 */
[
    uuid(0a781618-7e19-4a2c-8ec1-cf28db24247b),
    version(0.1.0)
]
interface IShortBuffer
{
    AsReadOnlyBuffer(
        [out] IShortBuffer** buffer);

    Compact();

    Duplicate(
        [out] IShortBuffer** buffer);

    Get(
        [out] Short* s);

    Get(
        [in] Integer index,
        [out] Short* s);

    Get(
        [out] Array<Short> dst);

    Get(
        [out] Array<Short> dst,
        [in] Integer offset,
        [in] Integer length);

    GetOrder(
        [out] IByteOrder** bo);

    HasArray(
        [out] Boolean* result);

    Put(
        [in] Short s);

    Put(
        [in] Integer index,
        [in] Short s);

    Put(
        [in] Array<Short> src);

    Put(
        [in] Array<Short> src,
        [in] Integer offset,
        [in] Integer length);

    Put(
        [in] IShortBuffer* src);

    Slice(
        [out] IShortBuffer** buffer);
}

}
}
