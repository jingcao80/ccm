//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace text {

/*
 * @Involve interface como::io::ISerializable
 * @Involve interface como::core::ICloneable
 */
[
    uuid(b2e89609-5020-4f1a-ae3b-3406c4021da1),
    version(0.1.0)
]
interface IDateFormatSymbols
{
    GetAmPmStrings(
        [out, callee] Array<String>* ampm);

    GetEras(
        [out, callee] Array<String>* eras);

    GetLocalPatternChars(
        [out] String* localPatternChars);

    GetMonths(
        [out, callee] Array<String>* months);

    GetShortMonths(
        [out, callee] Array<String>* months);

    GetShortWeekdays(
        [out, callee] Array<String>* weekdays);

    GetWeekdays(
        [out, callee] Array<String>* weekdays);

    GetZoneStrings(
        [out, callee] Array<Array<String>>* zoneStrings);

    SetAmPmStrings(
        [in] Array<String> newAmpms);

    SetEras(
        [in] Array<String> newEras);

    SetLocalPatternChars(
        [in] String newLocalPatternChars);

    SetMonths(
        [in] Array<String> newMonths);

    SetShortMonths(
        [in] Array<String> newShortMonths);

    SetShortWeekdays(
        [in] Array<String> newShortWeekdays);

    SetWeekdays(
        [in] Array<String> newWeekdays);

    SetZoneStrings(
        [in] Array<Array<String>> newZoneStrings);
}

}
}
