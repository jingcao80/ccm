//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace core {

interface ICharSequence;

[
    uuid(46d6e833-cb8a-4b12-9e3c-bfc25bf7c8f7),
    version(0.1.0)
]
interface IAppendable
{
    Append(
        [in] ICharSequence* csq);

    Append(
        [in] ICharSequence* csq,
        [in] Integer start,
        [in] Integer end);

    Append(
        [in] Char c);
}

}
}
