//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ISatellite.cdl"

namespace Universe {
namespace MilkyWay {
namespace SolarSystem {

[
    uuid(b1a08a58-761c-4c4c-81f2-ec7d71fcfdb3),
    version(0.1.0)
]
interface IMoon : ISatellite
{
    const String AROUND_PLANT_NAME = "Earth";
}

} // namespace SolarSystem
} // namespace MilkyWay
} // namespace Universe
