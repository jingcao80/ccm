//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::core::ICharSequence;
interface ccm::io::IByteBuffer;
interface ccm::io::ICharBuffer;
interface ccm::io::charset::ICodingErrorAction;
interface ccm::io::charset::ICoderResult;

namespace ccm {
namespace io {
namespace charset {

[
    uuid(1b6e3b85-c728-4a3f-a840-1d7b0eacc764),
    version(0.1.0)
]
interface ICharsetEncoder
{
    CanEncode(
        [in] Char c,
        [out] Boolean* result);

    CanEncode(
        [in] ICharSequence* cs,
        [out] Boolean* result);

    Encode(
        [in] ICharBuffer* cb,
        [out] IByteBuffer** bb);

    Encode(
        [in] ICharBuffer* cb,
        [out] IByteBuffer* bb,
        [in] Boolean endOfInput,
        [out] ICoderResult** result);

    Flush(
        [out] IByteBuffer* bb,
        [out] ICoderResult** result);

    GetAverageBytesPerChar(
        [out] Float* averageBytesPerChar);

    GetCharset(
        [out] ICharset** cs);

    GetMalformedInputAction(
        [out] ICodingErrorAction** action);

    GetMaxBytesPerChar(
        [out] Float* maxBytesPerChar);

    GetReplacement(
        [out, callee] Array<Byte>* replacement);

    GetUnmappableCharacterAction(
        [out] ICodingErrorAction** action);

    IsLegalReplacement(
        [in] Array<Byte> repl,
        [out] Boolean* isLegal);

    OnMalformedInput(
        [in] ICodingErrorAction* newAction);

    OnUnmappableCharacter(
        [in] ICodingErrorAction* newAction);

    ReplaceWith(
        [in] Array<Byte> newReplacement);

    Reset();
}

}
}
}
