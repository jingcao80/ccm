//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::text::IFormatField;
interface como::text::IFormatFieldDelegate;

namespace como {
namespace text {

[
    uuid(a847451b-46f3-441e-ba9f-ed0b37e5ebfa),
    version(0.1.0)
]
interface IFieldPosition
{
    GetBeginIndex(
        [out] Integer* index);

    GetEndIndex(
        [out] Integer* index);

    GetField(
        [out] Integer* field);

    GetFieldAttribute(
        [out] IFormatField** attribute);

    GetFieldDelegate(
        [out] IFormatFieldDelegate** delegate);

    SetBeginIndex(
        [in] Integer index);

    SetEndIndex(
        [in] Integer index);
}

}
}
