//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::util::IMapEntry;
interface como::util::INavigableSet;
interface como::util::ISortedMap;

namespace como {
namespace util {

/*
 * @Involve interface como::util::ISortedMap
 * @Involve interface como::util::IMap
 */
[
    uuid(db174312-1174-4777-8e66-e6f72359d0b8),
    version(0.1.0)
]
interface INavigableMap
{
    CeilingEntry(
        [in] IInterface* key,
        [out] IMapEntry&& entry);

    CeilingKey(
        [in] IInterface* key,
        [out] IInterface&& ceilingkey);

    DescendingKeySet(
        [out] INavigableSet&& keyset);

    DescendingMap(
        [out] INavigableMap&& map);

    FirstEntry(
        [out] IMapEntry&& entry);

    FloorEntry(
        [in] IInterface* key,
        [out] IMapEntry&& entry);

    FloorKey(
        [in] IInterface* key,
        [out] IInterface&& floorkey);

    HeadMap(
        [in] IInterface* toKey,
        [out] ISortedMap&& headmap);

    HeadMap(
        [in] IInterface* key,
        [in] Boolean inclusive,
        [out] INavigableMap&& headmap);

    HigherEntry(
        [in] IInterface* key,
        [out] IMapEntry&& entry);

    HigherKey(
        [in] IInterface* key,
        [out] IInterface&& higherkey);

    LastEntry(
        [out] IMapEntry&& entry);

    LowerEntry(
        [in] IInterface* key,
        [out] IMapEntry&& entry);

    LowerKey(
        [in] IInterface* key,
        [out] IInterface&& lowerkey);

    NavigableKeySet(
        [out] INavigableSet&& keyset);

    PollFirstEntry(
        [out] IMapEntry&& entry);

    PollLastEntry(
        [out] IMapEntry&& entry);

    SubMap(
        [in] IInterface* fromKey,
        [in] IInterface* toKey,
        [out] ISortedMap&& submap);

    SubMap(
        [in] IInterface* fromKey,
        [in] Boolean fromInclusive,
        [in] IInterface* toKey,
        [in] Boolean toInclusive,
        [out] INavigableMap&& submap);

    TailMap(
        [in] IInterface* fromKey,
        [out] ISortedMap&& tailmap);

    TailMap(
        [in] IInterface* fromKey,
        [in] Boolean inclusive,
        [out] INavigableMap&& tailmap);
}

}
}
