//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::io::IInputStream;
interface como::io::IOutputStream;
interface como::io::IPrintStream;
interface como::io::IPrintWriter;
interface como::io::IReader;
interface como::io::IWriter;

namespace como {
namespace util {

interface IEnumeration;
interface ISet;

/*
 * @Involve interface como::util::IHashtable;
 * @Involve interface como::util::IDictionary;
 * @Involve interface como::util::IMap;
 * @Involve interface como::core::ICloneable;
 * @Involve interface como::io::ISerializable;
 */
[
    uuid(417c6542-16e1-4542-b387-3f5075d73bee),
    version(0.1.0)
]
interface IProperties
{
    GetProperty(
        [in] String key,
        [out] String* value);

    GetProperty(
        [in] String key,
        [in] String defaultValue,
        [out] String* value);

    List(
        [in] IPrintStream* outstream);

    List(
        [in] IPrintWriter* outwriter);

    Load(
        [in] IInputStream* instream);

    Load(
        [in] IReader* reader);

    LoadFromXML(
        [in] IInputStream* instream);

    PropertyNames(
        [out] IEnumeration** names);

    Save(
        [in] IOutputStream* outstream,
        [in] String comments);

    SetProperty(
        [in] String key,
        [in] String value,
        [out] String* prevValue = nullptr);

    StringPropertyNames(
        [out] ISet&& names);

    Store(
        [in] IOutputStream* outstream,
        [in] String comment);

    Store(
        [in] IWriter* writer,
        [in] String comment);

    StoreToXML(
        [in] IOutputStream* os,
        [in] String comment);

    StoreToXML(
        [in] IOutputStream* os,
        [in] String comment,
        [in] String encoding);
}

}
}
