//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {

interface ICollection;
interface IIterator;
interface IList;
interface IListIterator;

/*
 * @Involve interface como::util::IList
 * @Involve interface como::util::ICollection
 * @Involve interface como::util::IRandomAccess
 * @Involve interface como::core::ICloneable
 * @Involve interface como::core::IIterable
 * @Involve interface como::io::ISerializable
 */
[
    uuid(d0dcbefa-d6ac-4f0e-96b7-e7697606f877),
    version(0.1.0)
]
interface IArrayList
{
    Add(
        [in] IInterface* obj,
        [out] Boolean* result = nullptr);

    Add(
        [in] Integer index,
        [in] IInterface* obj);

    AddAll(
        [in] ICollection* c,
        [out] Boolean* result = nullptr);

    AddAll(
        [in] Integer index,
        [in] ICollection* c,
        [out] Boolean* result = nullptr);

    Clear();

    Contains(
        [in] IInterface* obj,
        [out] Boolean& result);

    ContainsAll(
        [in] ICollection* c,
        [out] Boolean& result);

    EnsureCapacity(
        [in] Integer minCapacity);

    Equals(
        [in] IInterface* obj,
        [out] Boolean& result);

    Get(
        [in] Integer index,
        [out] IInterface&& obj);

    GetHashCode(
        [out] Integer& hash);

    GetIterator(
        [out] IIterator&& it);

    GetListIterator(
        [out] IListIterator&& it);

    GetListIterator(
        [in] Integer index,
        [out] IListIterator&& it);

    GetSize(
        [out] Integer& size);

    IndexOf(
        [in] IInterface* obj,
        [out] Integer& index);

    IsEmpty(
        [out] Boolean& empty);

    LastIndexOf(
        [in] IInterface* obj,
        [out] Integer& index);

    Remove(
        [in] IInterface* obj,
        [out] Boolean* result = nullptr);

    Remove(
        [in] Integer index,
        [out] IInterface** obj = nullptr);

    RemoveAll(
        [in] ICollection* c,
        [out] Boolean* result = nullptr);

    RetainAll(
        [in] ICollection* c,
        [out] Boolean* result = nullptr);

    Set(
        [in] Integer index,
        [in] IInterface* obj,
        [out] IInterface** prevObj = nullptr);

    SubList(
        [in] Integer fromIndex,
        [in] Integer toIndex,
        [out] IList&& subList);

    ToArray(
        [out, callee] Array<IInterface*>* objs);

    ToArray(
        [in] InterfaceID iid,
        [out, callee] Array<IInterface*>* objs);

    TrimToSize();
}

}
}
