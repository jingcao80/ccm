//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

/**
 * This file contains the definition of interface IPlanet.
 * IPlanet is an ICelestialBody which kind is planet.
 */

include "ICelestialBody.cdl"
include "ISatellite.cdl"

interface Universe.IStar;

namespace Universe {

[
    uuid(6fbd4882-ca56-4f46-8a9e-2efaff3c0528),
    version(0.1.0),
    description("This is the definition of IPlanet.")
]
interface IPlanet : ICelestialBody
{
    const CelestialBodyKind = planet;

    GetAroundStar(
        [out] IStar** star);

    GetDistanceToStar(
        [out] Double* distance);

    GetOrbitalPeriod(
        [out] Integer* hours);

    HasSatellite(
        [out] Boolean* hasSatellite);

    GetSatelliteNumber(
        [out] Integer* number);

    GetAllSatellites(
        [out] Array<ISatellite*>* satellites);

    GetAllSatellites(
        [out, callee] Array<ISatellite*>** satellites);
}

}  // namespace Universe
