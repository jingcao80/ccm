//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::util::IDate;

namespace ccm {
namespace util {

/*
 * @Involve interface ccm::util::ICalendar
 * @Involve interface ccm::io::ISerializable
 * @Involve interface ccm::core::ICloneable
 * @Involve interface ccm::core::IComparable
 */
[
    uuid(d6e54cfc-072f-4dba-98c3-b73d0931a53b),
    version(0.1.0)
]
interface IGregorianCalendar
{
    const Integer BC = 0;

    const Integer AD = 1;

    SetGregorianChange(
        [in] IDate* date);
}

}
}
