//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface libcore::io::IBufferIterator;

namespace libcore {
namespace util {

/*
 * @Involve interface ccm::util::ITimeZone
 * @Involve interface ccm::io::ISerializable
 * @Involve interface ccm::core::ICloneable
 */
[
    uuid(b06cc99d-8828-4e83-bb05-3ab04ac4b77b),
    version(0.1.0)
]
interface IZoneInfo
{
    FindTransitionIndex(
        [in] Long seconds,
        [out] Integer* index);

    GetOffsetsByUtcTime(
        [in] Long utcTimeInMillis,
        [out] Array<Integer> offsets,
        [out] Integer* total = nullptr);
}

[
    uuid(0b21624c-3400-44e0-84bc-d44dea940c9b),
    version(0.1.0)
]
interface IZoneInfoWallTime
{
    GetGmtOffset(
        [out] Integer* gmtoff);

    GetHour(
        [out] Integer* hour);

    GetIsDst(
        [out] Integer* isDst);

    GetMinute(
        [out] Integer* minute);

    GetMonth(
        [out] Integer* month);

    GetMonthDay(
        [out] Integer* monthDay);

    GetSecond(
        [out] Integer* second);

    GetWeekDay(
        [out] Integer* weekDay);

    GetYear(
        [out] Integer* year);

    GetYearDay(
        [out] Integer* yearDay);

    Localtime(
        [in] Integer timeSeconds,
        [in] IZoneInfo* zoneInfo);

    Mktime(
        [in] IZoneInfo* zoneInfo,
        [out] Integer* time);

    SetGmtOffset(
        [in] Integer gmtoff);

    SetHour(
        [in] Integer hour);

    SetIsDst(
        [in] Integer isDst);

    SetMinute(
        [in] Integer minute);

    SetMonth(
        [in] Integer month);

    SetMonthDay(
        [in] Integer monthDay);

    SetSecond(
        [in] Integer second);

    SetWeekDay(
        [in] Integer weekDay);

    SetYear(
        [in] Integer year);

    SetYearDay(
        [in] Integer yearDay);
}

}
}
