//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "libcore/io/IBufferIterator.cdl"
include "libcore/io/IIoBridge.cdl"
include "libcore/io/ILibcore.cdl"
include "libcore/io/IMemoryMappedFile.cdl"
include "libcore/io/IOs.cdl"

interface como::core::IAutoCloseable;

namespace libcore {
namespace io {

[
    uuid(cfaed610-0e3c-4e2a-a533-2fccc50ae541),
    version(0.1.0)
]
coclass CLibcore
{
    interface ILibcore;
}

[
    uuid(4fd4ee55-6fc3-4dd2-af89-e1a560cf707c),
    version(0.1.0)
]
coclass CMemoryMappedFile
{
    Constructor(
        [in] HANDLE address,
        [in] Long size);

    interface IMemoryMappedFile;
    interface IAutoCloseable;
}

}
}
