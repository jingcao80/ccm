//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace pisces {
namespace system {

[
    uuid(c5e4c12c-e52d-44d5-bbb3-55fda2d9eea8),
    version(0.1.0)
]
interface IStructStat
{
    /** Time of last access. */
    GetAtime(
        [out] Long* atime);

    /**
     * A file system-specific preferred I/O block size for this object.
     * For some file system types, this may vary from file to file.
     */
    GetBlksize(
        [out] Long* blksize);

    /** Number of blocks allocated for this object. */
    GetBlocks(
        [out] Long* blocks);

    /** Time of last status change. */
    GetCtime(
        [out] Long* ctime);

    /** Device ID of device containing file. */
    GetDev(
        [out] Long* dev);

    /** Group ID of file. */
    GetGid(
        [out] Integer* gid);

    /** File serial number (inode). */
    GetIno(
        [out] Long* ino);

    /** Mode (permissions) of file. */
    GetMode(
        [out] Integer* mode);

    /** Time of last data modification. */
    GetMtime(
        [out] Long* mtime);

    /** Number of hard links to the file. */
    GetNlink(
        [out] Long* nlink);

    /** Device ID (if file is character or block special). */
    GetRdev(
        [out] Long* rdev);

    /**
     * For regular files, the file size in bytes.
     * For symbolic links, the length in bytes of the pathname contained in the symbolic link.
     * For a shared memory object, the length in bytes.
     * For a typed memory object, the length in bytes.
     * For other file types, the use of this field is unspecified.
     */
    GetSize(
        [out] Long* size);

    /** User ID of file. */
    GetUid(
        [out] Integer* uid);
}

}
}
