//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace io {

[
    uuid(1a03d7ff-b6c9-4cb2-a30a-af6a5c6733e2),
    version(0.1.0)
]
interface IFileDescriptor
{
    GetInt(
        [out] Integer* fd);

    IsSocket(
        [out] Boolean* socket);

    SetInt(
        [in] Integer fd);

    Sync();

    Valid(
        [out] Boolean valid);
}

}
}
