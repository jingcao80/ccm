//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "comort/system/IBlockGuard.cdl"
include "comort/system/ICloseGuard.cdl"
include "comort/system/ISocketTagger.cdl"

interface como::IClassLoader;

namespace comort {
namespace system {

[
    uuid(dfa48353-9f1b-453d-a227-00f2390abe44),
    version(0.1.0)
]
coclass CPathClassLoader
{
    Constructor (
        [in] String classPath,
        [in] IClassLoader* parent);

    interface IClassLoader;
}

}
}
