//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface libcore::util::IZoneInfo;

namespace libcore {
namespace util {

[
    uuid(c2f5daa8-9f22-480b-8c63-fb9e79b7719b),
    version(0.1.0)
]
interface IZoneInfoDB
{}

[
    uuid(0ab77469-0ac6-4ced-bbc2-2c7eb0478a0e),
    version(0.1.0)
]
interface IZoneInfoDBTzData
{
    MakeTimeZone(
        [in] String id,
        [out] IZoneInfo** zone);
}

}
}
