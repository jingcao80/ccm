//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::io::IFileDescriptor;
interface como::net::IDatagramSocket;
interface como::net::ISocket;

namespace comort {
namespace system {

[
    uuid(bcf86319-3e1c-4c50-93cd-daea5797f296),
    version(0.1.0)
]
interface ISocketTagger
{
    Tag(
        [in] IFileDescriptor* socketDescriptor);

    Tag(
        [in] IDatagramSocket* socket);

    Tag(
        [in] ISocket* socket);

    Untag(
        [in] IFileDescriptor* socketDescriptor);

    Untag(
        [in] IDatagramSocket* socket);

    Untag(
        [in] ISocket* socket);
}

}
}
