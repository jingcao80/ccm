//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::core::IStackTraceElement;
interface ccm::io::IPrintStream;
interface ccm::io::IPrintWriter;

namespace ccm {
namespace core {

[
    uuid(b03ae37d-1d06-4a25-8d44-9790d292c9bf),
    version(0.1.0)
]
interface IStackTrace
{
    FillInStackTrace();

    GetStackTrace(
        [out, callee] Array<IStackTraceElement*>* stack);

    PrintStackTrace();

    PrintStackTrace(
        [in] IPrintStream* s);

    PrintStackTrace(
        [in] IPrintWriter* s);
}

}
}
