//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ccm/math/IBigDecimal.cdl"
include "ccm/math/IBigInteger.cdl"
include "ccm/math/IMathContext.cdl"
include "ccm/math/RoundingMode.cdl"

interface ccm::core::IComparable;
interface ccm::core::INumber;
interface ccm::io::ISerializable;
interface ccm::util::IRandom;

namespace ccm {
namespace math {

[
    uuid(c0f44da4-575b-44e6-b234-2208a28582ae),
    version(0.1.0)
]
coclass CBigDecimal
{
    Constructor(
        [in] Array<Char> arr,
        [in] Integer offset,
        [in] Integer len);

    Constructor(
        [in] Array<Char> arr,
        [in] Integer offset,
        [in] Integer len,
        [in] IMathContext* mc);

    Constructor(
        [in] Array<Char> arr);

    Constructor(
        [in] Array<Char> arr,
        [in] IMathContext* mc);

    Constructor(
        [in] String value);

    Constructor(
        [in] String value,
        [in] IMathContext* mc);

    Constructor(
        [in] Double value);

    Constructor(
        [in] Double value,
        [in] IMathContext* mc);

    Constructor(
        [in] IBigInteger* value);

    Constructor(
        [in] IBigInteger* value,
        [in] IMathContext* mc);

    Constructor(
        [in] IBigInteger* unscaledValue,
        [in] Integer scale);

    Constructor(
        [in] IBigInteger* unscaledValue,
        [in] Integer scale,
        [in] IMathContext* mc);

    Constructor(
        [in] Integer value);

    Constructor(
        [in] Integer value,
        [in] IMathContext* mc);

    Constructor(
        [in] Long value);

    Constructor(
        [in] Long value,
        [in] IMathContext* mc);

    interface IBigDecimal;
    interface INumber;
    interface IComparable;
    interface ISerializable;
}

[
    uuid(7a1ab981-ac06-4343-9746-db146876d3ac),
    version(0.1.0)
]
coclass CBigInteger
{
    Constructor(
        [in] Integer numBits,
        [in] IRandom* random);

    Constructor(
        [in] Integer bitLength,
        [in] Integer certainty,
        [in] IRandom* random);

    Constructor(
        [in] String value);

    Constructor(
        [in] String value,
        [in] Integer radix);

    Constructor(
        [in] Integer signum,
        [in] Array<Byte> magnitude);

    Constructor(
        [in] Array<Byte> value);

    interface IBigInteger;
    interface INumber;
    interface IComparable;
    interface ISerializable;
}

[
    uuid(3d32adb7-698c-4d2e-8421-fa2df3e0211c),
    version(0.1.0)
]
coclass CBigIntegerFactory
{
    interface IBigIntegerFactory;
}

[
    uuid(5542bfb6-c4d8-4fb2-a9b9-9683c61ad170),
    version(0.1.0)
]
coclass CMathContext
{
    Constructor(
        [in] Integer precision);

    Constructor(
        [in] Integer precision,
        [in] RoundingMode roundingMode);

    Constructor(
        [in] String s);

    interface IMathContext;
    interface ISerializable;
}

}
}
