//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "IStar.cdl"

namespace Universe {
namespace MilkyWay {
namespace SolarSystem {

[
    uuid(03b13c47-0982-46ba-bbbe-f43557df6ec9),
    version(0.1.0)
]
interface ISun : IStar
{
    GetDistanceToEarth(
        [out] Double* distance);
}

} // namespace SolarSystem
} // namespace MilkyWay
} // namespace Universe
