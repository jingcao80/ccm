//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

[
    uuid(f0a35bbc-25aa-4156-99f1-fa6e01bd8255),
    uri("http://como.org/component/test/ReferenceTypeTest.so")
]
module ReferenceTypeTest
{

namespace como {
namespace test {

[
    uuid(b2a278ee-f571-415e-bfaa-e8b305be3c65),
    version(0.1.0)
]
interface IFoo
{
    Foo(
        [in] Integer value,
        [out] Integer& result);
}

[
    uuid(beb8cc88-4a4f-4d97-9520-b6f4fe89ec10),
    version(0.1.0)
]
interface IBar
{
    Bar(
        [in] String name,
        [out] String& id);
}

[
    uuid(6103fa48-3f22-4769-acef-688a7d5a0590),
    version(0.1.0)
]
interface IFooBar
{
    FooBar(
        [in] IFoo* foo,
        [out] IBar&& bar);
}

[
    uuid(c39abf6b-4daf-4572-be0f-962a6a7b8639),
    version(0.1.0)
]
coclass CFooBar
{
    Constructor(
        [in] Integer initValue);

    interface IFoo;
    interface IBar;
    interface IFooBar;
}

} // namespace test
} // namespace como

}
