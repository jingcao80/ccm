//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {
namespace concurrent {
namespace atomic {

/*
 * @Involve interface ccm:core::INumber
 * @Involve interface ccm::io::ISerializable
 */
[
    uuid(991e8db3-d281-4acc-926b-ad1b1e3e2688),
    version(0.1.0)
]
interface IAtomicLong
{
    AddAndGet(
        [in] Long delta,
        [out] Long* value);

    CompareAndSet(
        [in] Long expect,
        [in] Long update,
        [out] Boolean* succeeded = nullptr);

    DecrementAndGet(
        [out] Long* value);

    Get(
        [out] Long* value);

    GetAndAdd(
        [in] Long delta,
        [out] Long* prevValue);

    GetAndDecrement(
        [out] Long* prevValue);

    GetAndIncrement(
        [out] Long* prevValue);

    GetAndSet(
        [in] Long newValue,
        [out] Long* prevValue);

    IncrementAndGet(
        [out] Long* value);

    LzaySet(
        [in] Long value);

    Set(
        [in] Long value);

    WeakCompareAndSet(
        [in] Long expect,
        [in] Long update,
        [out] Boolean* succeeded = nullptr);
}

}
}
}
}
