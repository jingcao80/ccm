//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::security::IProvider;

namespace ccm {
namespace security {

/*
 * @Involve interface ccm::util::IRandom
 * @Involve interface ccm::io:ISerializable
 */
[
    uuid(a9d0a2ef-0248-448d-ae16-2ff4df8ab0d7),
    version(0.1.0)
]
interface ISecureRandom
{
    GenerateSeed(
        [in] Integer numBytes,
        [out, callee] Array<Byte>* seed);

    GetAlgorithm(
        [out] String* algorithm);

    GetProvider(
        [out] IProvider** provider);

    SetSeed(
        [in] Array<Byte> seed);
}

}
}
