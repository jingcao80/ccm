//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

[
    uuid(3657416d-4638-4843-a0b9-eb7ef1794495),
    url("http://ccm.org/component/library/libcore.so")
]
module libcore
{

include "ccm/core.cdl"
include "ccm/io.cdl"
include "ccm/core2.cdl"
include "ccm/util.cdl"
include "ccmrt/system.cdl"

}
