//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace io {

/*
 * @involve ccm::io::ICloseable
 * @involve ccm::core::IAutoCloseable
 */
[
    uuid(ffea83b0-bb5d-4a13-b9e8-9a430b97e854),
    version(0.1.0)
]
interface IInputStream
{
    Available(
        [out] Integer* number);

    Close();

    IsMarkSupported(
        [out] Boolean* supported);

    Mark(
        [in] Integer readLimit);

    Read(
        [out] Integer* value);

    Read(
        [in] Array<Byte> buffer,
        [out] Integer* number);

    Read(
        [in] Array<Byte> buffer,
        [in] Integer offset,
        [in] Integer size,
        [out] Integer* number);

    Reset();

    Skip(
        [in] Long byteCount,
        [out] Long* number);
}

}
}
