//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::util::IComparator;

namespace como {
namespace util {

/*
 * @Involve interface como::util::ISet
 * @Involve interface como::util::ICollection
 * @Involve interface como::core::IIterable
 */
[
    uuid(87972ee6-547a-4ae5-b17d-a7e8f8ec794a),
    version(0.1.0)
]
interface ISortedSet
{
    Add(
        [in] IInterface* obj,
        [out] Boolean* modified = nullptr);

    Comparator(
        [out] IComparator&& comparator);

    First(
        [out] IInterface&& element);

    GetIterator(
        [out] IIterator&& it);

    HeadSet(
        [in] IInterface* toElement,
        [out] ISortedSet&& headset);

    Last(
        [out] IInterface&& element);

    SubSet(
        [in] IInterface* fromElement,
        [in] IInterface* toElement,
        [out] ISortedSet&& subset);

    TailSet(
        [in] IInterface* fromElement,
        [out] ISortedSet&& tailset);
}

}
}
