//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::util::ITimeZone;
interface ccm::util::calendar::ICalendarDate;
interface ccm::util::calendar::IEra;

namespace ccm {
namespace util {
namespace calendar {

[
    uuid(203ce39d-2cb3-45ec-a618-5f674a2494b8),
    version(0.1.0)
]
interface ICalendarSystem
{
    GetEra(
        [in] String eraName,
        [out] IEra** era);

    GetEras(
        [out, callee] Array<IEra*>* eras);

    GetCalendarDate(
        [out] ICalendarDate** date);

    GetCalendarDate(
        [in] Long millis,
        [out] ICalendarDate** date);

    GetCalendarDate(
        [in] Long millis,
        [in] ICalendarDate* inDate,
        [out] ICalendarDate** outDate);

    GetCalendarDate(
        [in] Long millis,
        [in] ITimeZone* zone,
        [out] ICalendarDate** date);

    GetMonthLength(
        [in] ICalendarDate* date,
        [out] Integer months);

    GetName(
        [out] String* name);

    GetNthDayOfWeek(
        [in] Integer nth,
        [in] Integer dayOfWeek,
        [in] ICalendarDate* inDate,
        [out] ICalendarDate** outDate);

    GetTime(
        [in] ICalendarDate* date,
        [out] Long* time);

    GetWeekLength(
        [out] Integer* weeks);

    GetYearLength(
        [in] ICalendarDate* date,
        [out] Integer* years);

    GetYearLengthInMonths(
        [in] ICalendarDate* date,
        [out] Integer* years);

    NewCalendarDate(
        [out] ICalendarDate** date);

    NewCalendarDate(
        [in] ITimeZone* zone,
        [out] ICalendarDate** date);

    Normalize(
        [in] ICalendarDate* date,
        [out] Boolean* result);

    SetEra(
        [in] ICalendarDate* date,
        [in] String eraName);

    SetTimeOfDay(
        [in] ICalendarDate* date,
        [in] Integer timeOfDay);

    Validate(
        [in] ICalendarDate* date,
        [out] Boolean* result);
}

}
}
}
