//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::util::IList;

namespace como {
namespace util {
namespace locale {

[
    uuid(527ad6e7-ef79-4133-8fc1-a38b614827ba),
    version(0.1.0)
]
interface ILanguageTag
{
    const String PRIVATEUSE = "x";

    const String PRIVUSE_VARIANT_PREFIX = "lvariant";

    const String SEP = "-";

    const String UNDETERMINED = "und";

    GetExtensions(
        [out] IList** extensions);

    GetExtlangs(
        [out] IList** extlangs);

    GetLanguage(
        [out] String* language);

    GetPrivateuse(
        [out] String* privateuse);

    GetRegion(
        [out] String* region);

    GetScript(
        [out] String* script);

    GetVariants(
        [out] IList** variants);
}

}
}
}
