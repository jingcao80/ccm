//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::core::IThread;

namespace ccm {
namespace core {

[
    uuid(22b24f1e-45ec-4669-86c8-a75cd6af7e2a),
    version(0.1.0)
]
interface IRuntime
{
    AddShutdownHook(
        [in] IThread* hook);

    AvailableProcessors(
        [out] Integer* ncpu);

    Exit(
        [in] Integer status);
}

[
    uuid(70d502ac-f307-4b5b-9b36-afe7ee687b7b),
    version(0.1.0)
]
interface IRuntimeFactory
{
    GetRuntime(
        [out] IRuntime** runtime);
}

}
}
