//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::io::ISerializable;

namespace ccm {
namespace core {

[
    uuid(df471c09-381f-40c4-9e24-c92b31dd9146),
    version(0.1.0)
]
coclass CBoolean
{
    constructor(
           [in] Boolean value);

   interface IBoolean;
   interface ISerializable;
   interface IComparable;
}

[
    uuid(bdf665c0-8a7a-4621-ba55-e6a097dfc85d),
    version(0.1.0)
]
coclass CByte
{
    constructor(
        [in] Byte value);

    interface IByte;
    interface INumber;
    interface ISerializable;
    interface IComparable;
}

[
    uuid(10e6419e-b8d0-44be-b309-54086eb3e560),
    version(0.1.0)
]
coclass CString
{
    constructor(
        [in] String str);

    interface ISerializable;
    interface ICharSequence;
    interface IComparable;
    interface IString;
}

[
    uuid(8c3a55f1-63c5-4abd-b68c-46773877a655),
    version(0.1.0)
]
coclass CStringBuffer
{
    constructor();

    constructor(
        [in] Integer capacity);

    constructor(
        [in] String str);

    constructor(
        [in] ICharSequence* seq);

    interface ISerializable;
    interface ICharSequence;
    interface IStringBuffer;
}

[
    uuid(cbc6b55a-c06e-4ddc-b7f8-f0cc0bf94ff9),
    version(0.1.0)
]
coclass CStringBuilder
{
    constructor();

    constructor(
        [in] Integer capacity);

    constructor(
        [in] String str);

    constructor(
        [in] ICharSequence* seq);

    interface ISerializable;
    interface ICharSequence;
    interface IStringBuilder;
}

}
}
