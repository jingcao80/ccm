//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::core::IAppendable;

namespace como {
namespace misc {

[
    uuid(6bb0744f-9dfe-451c-a68b-3e2c3bde5aa3),
    version(0.1.0)
]
interface IFloatingDecimalBinaryToASCIIConverter
{
    AppendTo(
        [in] IAppendable* buf);

    DecimalDigitsExact(
        [out] Boolean& exact);

    DigitsRoundedUp(
        [out] Boolean& roundedUp);

    GetDecimalExponent(
        [out] Integer& exponent);

    GetDigits(
        [out] Array<Char>& digits,
        [out] Integer& number);

    IsExceptional(
        [out] Boolean& exceptional);

    IsNegative(
        [out] Boolean& neg);

    ToFormatString(
        [out] String& str);
}

[
    uuid(691e4ffb-5b88-40de-ae6e-12072672fbbc),
    version(0.1.0)
]
interface IFloatingDecimalASCIIToBinaryConverter
{
    DoubleValue(
        [out] Double& value);

    FloatValue(
        [out] Float& value);
}

}
}
