//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ccm/util/Exceptions.cdl"
include "ccm/util/IArrayList.cdl"
include "ccm/util/ICollection.cdl"
include "ccm/util/IDate.cdl"
include "ccm/util/IDictionary.cdl"
include "ccm/util/IEnumeration.cdl"
include "ccm/util/IHashtable.cdl"
include "ccm/util/IHashMap.cdl"
include "ccm/util/IHashSet.cdl"
include "ccm/util/IIterator.cdl"
include "ccm/util/ILinkedHashMap.cdl"
include "ccm/util/ILinkedHashSet.cdl"
include "ccm/util/IList.cdl"
include "ccm/util/IListIterator.cdl"
include "ccm/util/ILocale.cdl"
include "ccm/util/IMap.cdl"
include "ccm/util/IProperties.cdl"
include "ccm/util/IRandom.cdl"
include "ccm/util/IRandomAccess.cdl"
include "ccm/util/ISet.cdl"
include "ccm/util/IStringTokenizer.cdl"
include "ccm/util/ITimeZone.cdl"
include "ccm/util/calendar/IBaseCalendar.cdl"
include "ccm/util/calendar/ICalendarDate.cdl"
include "ccm/util/calendar/ICalendarSystem.cdl"
include "ccm/util/calendar/IEra.cdl"
include "ccm/util/calendar/IGregorian.cdl"
include "ccm/util/calendar/IJulianCalendar.cdl"
include "ccm/util/calendar/ILocalGregorianCalendar.cdl"
include "ccm/util/concurrent/IConcurrentMap.cdl"
include "ccm/util/concurrent/atomic/IAtomicInteger.cdl"
include "ccm/util/concurrent/atomic/IAtomicLong.cdl"
include "ccm/util/regex/Exceptions.cdl"
include "ccm/util/regex/IMatcher.cdl"
include "ccm/util/regex/IMatchResult.cdl"
include "ccm/util/regex/IPattern.cdl"

interface ccm::core::ICloneable;
interface ccm::core::IComparable;
interface ccm::core::IIterable;
interface ccm::core::INumber;
interface ccm::io::ISerializable;

namespace ccm {
namespace util {

[
    uuid(7dbd4e0a-4bf2-4ccb-a4e9-bfe232b40ba4),
    version(0.1.0)
]
coclass CArrayList
{
    Constructor();

    Constructor(
        [in] Integer initialCapacity);

    Constructor(
        [in] ICollection* c);

    interface IArrayList;
    interface IList;
    interface ICollection;
    interface IRandomAccess;
    interface IIterable;
    interface ICloneable;
    interface ISerializable;
}

[
    uuid(57b9bd7b-d0d5-42c5-9784-202614517a4f),
    version(0.1.0)
]
coclass CDate
{
    Constructor();

    Constructor(
        [in] Long date);

    Constructor(
        [in] Integer year,
        [in] Integer month,
        [in] Integer date);

    Constructor(
        [in] Integer year,
        [in] Integer month,
        [in] Integer date,
        [in] Integer hrs,
        [in] Integer min);

    Constructor(
        [in] Integer year,
        [in] Integer month,
        [in] Integer date,
        [in] Integer hrs,
        [in] Integer min,
        [in] Integer sec);

    Constructor(
        [in] String s);

    interface IDate;
    interface ICloneable;
    interface IComparable;
    interface ISerializable;
}

[
    uuid(afe87a5a-0e0b-4c33-975e-2ec5caa60afc),
    version(0.1.0)
]
coclass CHashMap
{
    Constructor();

    Constructor(
        [in] Integer initialCapacity);

    Constructor(
        [in] IMap* m);

    Constructor(
        [in] Integer initialCapacity,
        [in] Float loadFactor);

    interface IHashMap;
    interface IMap;
    interface ICloneable;
    interface ISerializable;
}

[
    uuid(3b1f6a9d-3d2b-43ab-b61f-caa766e84303),
    version(0.1.0)
]
coclass CHashSet
{
    Constructor();

    Constructor(
        [in] ICollection* c);

    Constructor(
        [in] Integer initialCapacity);

    Constructor(
        [in] Integer initialCapacity,
        [in] Float loadFactor);

    Constructor(
        [in] Integer initialCapacity,
        [in] Float loadFactor,
        [in] Boolean dummy);

    interface IHashSet;
    interface ISet;
    interface ICollection;
    interface IIterable;
    interface ISerializable;
    interface ICloneable;
}

[
    uuid(10c87f0c-91e6-4fa1-905e-8ce9f513318f),
    version(0.1.0)
]
coclass CHashtable
{
    Constructor();

    Constructor(
        [in] Integer initialCapacity);

    Constructor(
        [in] Integer initialCapacity,
        [in] Float loadFactor);

    Constructor(
        [in] IMap* t);

    interface IHashtable;
    interface IDictionary;
    interface IMap;
    interface ICloneable;
    interface ISerializable;
}

[
    uuid(737c1ff9-c4b3-4d55-a67f-160a411d289b),
    version(0.1.0)
]
coclass CLinkedHashMap
{
    Constructor();

    Constructor(
        [in] Integer initialCapacity);

    Constructor(
        [in] Integer initialCapacity,
        [in] Float loadFactor);

    Constructor(
        [in] Integer initialCapacity,
        [in] Float loadFactor,
        [in] Boolean accessOrder);

    Constructor(
        [in] IMap* m);

    interface ILinkedHashMap;
    interface IHashMap;
    interface IMap;
    interface ICloneable;
    interface ISerializable;
}

[
    uuid(2a5b0a37-7877-4ee5-9b3a-439538f70354),
    version(0.1.0)
]
coclass CLinkedHashSet
{
    Constructor();

    Constructor(
        [in] ICollection* c);

    Constructor(
        [in] Integer initialCapacity);

    Constructor(
        [in] Integer initialCapacity,
        [in] Float loadFactor);

    interface ILinkedHashSet;
    interface IHashSet;
    interface ISet;
    interface ICollection;
    interface IIterable;
    interface ISerializable;
    interface ICloneable;
}

[
    uuid(2f6a7390-6aed-4f7d-863e-3f007635ba14),
    version(0.1.0)
]
coclass CProperties
{
    Constructor();

    Constructor(
        [in] IProperties* defaults);

    interface IProperties;
    interface IHashtable;
    interface IDictionary;
    interface IMap;
    interface ICloneable;
    interface ISerializable;
}

[
    uuid(1d590d6f-70ee-497a-b8a9-e99212e04f53),
    version(0.1.0)
]
coclass CRandom
{
    Constructor();

    Constructor(
        [in] Long seed);

    interface IRandom;
    interface ISerializable;
}

[
    uuid(6858c0ba-e3a0-48fd-8f22-bbdc4503d83d),
    version(0.1.0)
]
coclass CStringTokenizer
{
    Constructor(
        [in] String str,
        [in] String delim,
        [in] Boolean returnDelims);

    Constructor(
        [in] String str,
        [in] String delim);

    Constructor(
        [in] String str);

    interface IStringTokenizer;
    interface IEnumeration;
}

namespace calendar {

[
    uuid(d8b9fb39-2e68-4209-8cd3-9a2f0235f9e2),
    version(0.1.0)
]
coclass CCalendarSystemFactory
{
    interface ICalendarSystemFactory;
}

[
    uuid(40eab8b9-84da-4399-a171-ce260a17204a),
    version(0.1.0)
]
coclass CEra
{
    Constructor(
        [in] String name,
        [in] String abbr,
        [in] Long since,
        [in] Boolean localTime);

    interface IEra;
}

[
    uuid(f726de31-d4f4-440b-b8a5-dfb25fea88d2),
    version(0.1.0)
]
coclass CGregorian
{
    // @hide
    Constructor();

    interface IGregorian;
    interface IBaseCalendar;
    interface ICalendarSystem;
}

[
    uuid(d6038b88-1454-4a8a-a17d-dbf16151a36b),
    version(0.1.0)
]
coclass CJulianCalendar
{
    // @hide
    Constructor();

    interface IJulianCalendar;
    interface IBaseCalendar;
    interface ICalendarSystem;
}

[
    uuid(4b4a5802-2e14-45cf-9894-2c9645972a5c),
    version(0.1.0)
]
coclass CLocalGregorianCalendar
{
    // @hide
    Constructor(
        [in] String name,
        [in] Array<IEra*> eras);

    interface ILocalGregorianCalendar;
    interface IBaseCalendar;
    interface ICalendarSystem;
}

}

namespace concurrent {

namespace atomic {

[
    uuid(37e94445-0ee6-460f-9105-4afed59d6586),
    version(0.1.0)
]
coclass CAtomicInteger
{
    Constructor();

    Constructor(
        [in] Integer initialValue);

    interface IAtomicInteger;
    interface INumber;
    interface ISerializable;
}

[
    uuid(067d7bcc-d79c-43be-ada6-459adf04619e),
    version(0.1.0)
]
coclass CAtomicLong
{
    Constructor();

    Constructor(
        [in] Long initialValue);

    interface IAtomicLong;
    interface INumber;
    interface ISerializable;
}

}

}

namespace regex {

[
    uuid(698f1b9a-dd5e-4ae4-924c-c1addd038571),
    version(0.1.0)
]
coclass CPatternFactory
{
    interface IPatternFactory;
}

}
}
}
