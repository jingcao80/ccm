//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace libcore {
namespace io {

[
    uuid(c76aba68-5070-4475-9dea-232106fa27ea),
    version(0.1.0)
]
interface IBufferIterator
{
    Pos(
        [out] Integer* offset);

    ReadByte(
        [out] Byte* result);

    ReadByteArray(
        [out] Array<Byte> dst,
        [in] Integer dstOffset,
        [in] Integer byteCount);

    ReadInteger(
        [out] Integer* result);

    ReadIntegerArray(
        [out] Array<Integer> dst,
        [in] Integer dstOffset,
        [in] Integer intCount);

    ReadShort(
        [out] Short* result);

    Seek(
        [in] Integer offset);

    Skip(
        [in] Integer byteCount);
}

}
}
