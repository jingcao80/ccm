//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace io {

/*
 * @Involve interface como::io::IBuffer;
 * @Involve interface como::core::IComparable;
 */
[
    uuid(e0f0ef95-b242-4716-bae7-d4e047fda555),
    version(0.1.0)
]
interface ILongBuffer
{
    AsReadOnlyBuffer(
        [out] ILongBuffer** buffer);

    Compact();

    Duplicate(
        [out] ILongBuffer** buffer);

    Get(
        [out] Long* l);

    Get(
        [in] Integer index,
        [out] Long* l);

    Get(
        [out] Array<Long> dst);

    Get(
        [out] Array<Long> dst,
        [in] Integer offset,
        [in] Integer length);

    GetOrder(
        [out] IByteOrder** bo);

    HasArray(
        [out] Boolean* result);

    Put(
        [in] Long l);

    Put(
        [in] Integer index,
        [in] Long l);

    Put(
        [in] Array<Long> src);

    Put(
        [in] Array<Long> src,
        [in] Integer offset,
        [in] Integer length);

    Put(
        [in] ILongBuffer* src);

    Slice(
        [out] ILongBuffer** buffer);
}

}
}
