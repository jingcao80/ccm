//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace jing {
namespace icu {
namespace text {

enum ITimeZoneNamesNameType
{
    /**
     * Long display name, such as "Eastern Time".
     */
    ONG_GENERIC,

    /**
     * Long display name for standard time, such as "Eastern Standard Time".
     */
    LONG_STANDARD,

    /**
     * Long display name for daylight saving time, such as "Eastern Daylight Time".
     */
    LONG_DAYLIGHT,

    /**
     * Short display name, such as "ET".
     */
    SHORT_GENERIC,

    /**
     * Short display name for standard time, such as "EST".
     */
    SHORT_STANDARD,

    /**
     * Short display name for daylight saving time, such as "EDT".
     */
    SHORT_DAYLIGHT,

    /**
     * Exemplar location name, such as "Los Angeles".
     */
    EXEMPLAR_LOCATION,
}

[
    uuid(b1f01233-3da2-4b26-a041-519317137cf7),
    version(0.1.0)
]
interface ITimeZoneNames
{

}

}
}
}
