//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "pisces/system/IStructAddrinfo.cdl"
include "pisces/system/IStructCapUserData.cdl"
include "pisces/system/IStructCapUserHeader.cdl"
include "pisces/system/IStructFlock.cdl"
include "pisces/system/IStructGroupReq.cdl"
include "pisces/system/IStructGroupSourceReq.cdl"
include "pisces/system/IStructIfaddrs.cdl"
include "pisces/system/IStructLinger.cdl"
include "pisces/system/IStructPasswd.cdl"
include "pisces/system/IStructPollfd.cdl"
include "pisces/system/IStructStat.cdl"
include "pisces/system/IStructStatVfs.cdl"
include "pisces/system/IStructTimeval.cdl"
include "pisces/system/IStructUcred.cdl"
include "pisces/system/IStructUtsname.cdl"
