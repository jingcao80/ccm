//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

const Integer ICONST1 = 1;

namespace como {
namespace test {

const Integer ICONST2 = 2;

namespace reflection {

const Integer ICONST3 = 3;

const Float FCONST = ICONST3;

const Double DCONST = FCONST;

}

}
}

const Byte BCONST = ICONST1 + 5;

const Char CCONST = BCONST;

const Short SCONST = CCONST * 10;
