//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace comort {
namespace system {

[
    uuid(17faccd7-40f0-43ba-a68a-b127bf175642),
    version(0.1.0)
]
interface IBlockGuardPolicy
{
    OnWriteToDisk();

    OnReadFromDisk();

    OnNetwork();

    OnUnbufferedIO();

    GetPolicyMask(
        [out] Integer* mask);
}

[
    uuid(eca31f7d-c4f5-4bb4-af3e-c015af278c29),
    version(0.1.0)
]
interface IBlockGuard
{
    const Integer DISALLOW_DISK_WRITE = 0x01;
    const Integer DISALLOW_DISK_READ = 0x02;
    const Integer DISALLOW_NETWORK = 0x04;
    const Integer PASS_RESTRICTIONS_VIA_RPC = 0x08;
    const Integer PENALTY_LOG = 0x10;
    const Integer PENALTY_DIALOG = 0x20;
    const Integer PENALTY_DEATH = 0x40;

    GetLaxPolicy(
        [out] IBlockGuardPolicy** policy);

    GetThreadPolicy(
        [out] IBlockGuardPolicy** policy);

    SetThreadPolicy(
        [in] IBlockGuardPolicy* policy);
}

}
}
