//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::IInterface;
interface ccm::io::IByteBuffer;
interface ccm::io::IFileDescriptor;
interface ccm::net::IDatagramPacket;
interface ccm::net::IInetAddress;
interface ccm::net::IInetSocketAddress;
interface libcore::io::IOs;

namespace libcore {
namespace io {

[
    uuid(e20a68e0-d3fa-4415-ba77-b6e663f1ac8c),
    version(0.1.0)
]
interface IoBridge
{
    Available(
        [in] IFileDescriptor* fd,
        [out] Integer* number);

    Bind(
        [in] IFileDescriptor* fd,
        [in] IInetAddress* address,
        [in] Integer port);

    Connect(
        [in] IFileDescriptor* fd,
        [in] IInetAddress* inetAddress,
        [in] Integer port);

    Connect(
        [in] IFileDescriptor* fd,
        [in] IInetAddress* inetAddress,
        [in] Integer port,
        [in] Integer timeoutMs);

    CloseAndSignalBlockedThreads(
        [in] IFileDescriptor* fd);

    IsConnected(
        [in] IFileDescriptor* fd,
        [in] IInetAddress* inetAddress,
        [in] Integer port,
        [in] Integer timeoutMs,
        [in] Integer remainingTimeoutMs,
        [out] Boolean connected);

    GetLocalInetSocketAddress(
        [in] IFileDescriptor* fd,
        [out] IInetSocketAddress** socket);

    GetSocketOption(
        [in] IFileDescriptor* fd,
        [in] Integer option,
        [out] IInterface** socket);

    Open(
        [in] String path,
        [in] Integer flags,
        [out] IFileDescriptor** fd);

    Poll(
        [in] IFileDescriptor* fd,
        [in] Integer events,
        [in] Integer timeout);

    Read(
        [in] IFileDescriptor* fd,
        [out] Array<Byte> bytes,
        [in] Integer byteOffset,
        [in] Integer byteCount,
        [out] Integer* number);

    Recvfrom(
        [in] Boolean isRead,
        [in] IFileDescriptor* fd,
        [out] Array<Byte> bytes,
        [in] Integer byteOffset,
        [in] Integer byteCount,
        [in] Integer flags,
        [in] IDatagramPacket* packet,
        [in] Boolean isConnected,
        [out] Integer* number);

    Recvfrom(
        [in] Boolean isRead,
        [in] IFileDescriptor* fd,
        [in] IByteBuffer* buffer,
        [in] Integer flags,
        [in] IDatagramPacket* packet,
        [in] Boolean isConnected,
        [out] Integer* number);

    Sendto(
        [in] IFileDescriptor* fd,
        [in] Array<Byte> bytes,
        [in] Integer byteOffset,
        [in] Integer byteCount,
        [in] Integer flags,
        [in] IInetAddress* inetAddress,
        [in] Integer port,
        [out] Integer* number);

    Sendto(
        [in] IFileDescriptor* fd,
        [in] IByteBuffer* buffer,
        [in] Integer flags,
        [in] IInetAddress* inetAddress,
        [in] Integer port,
        [out] Integer* number);

    SetSocketOption(
        [in] IFileDescriptor* fd,
        [in] Integer option,
        [in] IInterface* value);

    Socket(
        [in] Integer domain,
        [in] Integer type,
        [in] Integer protocol,
        [out] IFileDescriptor** fd);

    Write(
        [in] IFileDescriptor* fd,
        [in] Array<Byte> bytes,
        [in] Integer byteOffset,
        [in] Integer byteCount);
}

}
}
