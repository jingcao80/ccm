//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ccm/math/IBigDecimal.cdl"
include "ccm/math/IBigInteger.cdl"

interface ccm::core::IComparable;
interface ccm::core::INumber;
interface ccm::io::ISerializable;
interface ccm::util::IRandom;

namespace ccm {
namespace math {

[
    uuid(7a1ab981-ac06-4343-9746-db146876d3ac),
    version(0.1.0)
]
coclass CBigInteger
{
    Constructor(
        [in] Integer numBits,
        [in] IRandom* random);

    Constructor(
        [in] Integer bitLength,
        [in] Integer certainty,
        [in] IRandom* random);

    Constructor(
        [in] String value);

    Constructor(
        [in] String value,
        [in] Integer radix);

    Constructor(
        [in] Integer signum,
        [in] Array<Byte> magnitude);

    Constructor(
        [in] Array<Byte> value);

    interface IBigInteger;
    interface INumber;
    interface IComparable;
    interface ISerializable;
}

[
    uuid(3d32adb7-698c-4d2e-8421-fa2df3e0211c),
    version(0.1.0)
]
coclass CBigIntegerFactory
{
    interface IBigIntegerFactory;
}

}
}
