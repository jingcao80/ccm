//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {

interface ICollection;
interface IIterator;

/*
 * @Involve interface como::util::ICollection
 * @Involve interface como::core::IIterable
 */
[
    uuid(163ff32d-c566-4666-8b18-73b5062751c0),
    version(0.1.0)
]
interface ISet
{
    Add(
        [in] IInterface* obj,
        [out] Boolean* modified = nullptr);

    AddAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    Clear();

    Contains(
        [in] IInterface* obj,
        [out] Boolean* result);

    ContainsAll(
        [in] ICollection* c,
        [out] Boolean* result);

    Equals(
        [in] IInterface* obj,
        [out] Boolean& result);

    GetHashCode(
        [out] Integer& hash);

    GetIterator(
        [out] IIterator&& it);

    GetSize(
        [out] Integer* size);

    IsEmpty(
        [out] Boolean* result);

    Remove(
        [in] IInterface* obj,
        [out] Boolean* contained = nullptr);

    RemoveAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    RetainAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    ToArray(
        [out, callee] Array<IInterface*>* objs);

    ToArray(
        [in] InterfaceID iid,
        [out, callee] Array<IInterface*>* objs);
}

}
}
