//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::text::IAttributedCharacterIterator;
interface ccm::text::IAttributedCharacterIteratorAttribute;
interface ccm::util::IMap;

namespace ccm {
namespace text {

[
    uuid(b3004d6b-0223-4bcb-8b6d-7824de3aeb3a),
    version(0.1.0)
]
interface IAttributedString
{
    AddAttribute(
        [in] IAttributedCharacterIteratorAttribute* attribute,
        [in] IInterface* value);

    AddAttribute(
        [in] IAttributedCharacterIteratorAttribute* attribute,
        [in] IInterface* value,
        [in] Integer beginIndex,
        [in] Integer endIndex);

    AddAttributes(
        [in] IMap* attributes,
        [in] Integer beginIndex,
        [in] Integer endIndex);

    GetIterator(
        [out] IAttributedCharacterIterator** it);

    GetIterator(
        [in] Array<IAttributedCharacterIteratorAttribute*> attributes,
        [out] IAttributedCharacterIterator** it);

    GetIterator(
        [in] Array<IAttributedCharacterIteratorAttribute*> attributes,
        [in] Integer beginIndex,
        [in] Integer endIndex,
        [out] IAttributedCharacterIterator** it);
}

}
}
