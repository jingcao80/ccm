//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::core::ICharSequence;
interface ccm::core::IStringBuffer;

namespace ccm {
namespace util {
namespace regex {

interface IMatchResult;
interface IPattern;

[
    uuid(59e2bbf1-fc3a-4525-9eb0-cfa32d7c75c7),
    version(0.1.0)
]
interface IMatcher
{
    AppendReplacement(
        [in] IStringBuffer* sb,
        [in] String replacement);

    AppendTail(
        [in] IStringBuffer* sb);

    End(
        [out] Integer* index);

    End(
        [in] Integer group,
        [out] Integer* index);

    End(
        [in] String name,
        [out] Integer* index);

    Find(
        [out] Boolean* result);

    Find(
        [in] Integer start,
        [out] Boolean* result);

    Group(
        [out] String* subseq);

    Group(
        [in] Integer group,
        [out] String* subseq);

    Group(
        [in] String name,
        [out] String* subseq);

    GroupCount(
        [out] Integer* number);

    HasAnchoringBounds(
        [out] Boolean* result);

    HasTransparentBounds(
        [out] Boolean* result);

    HitEnd(
        [out] Boolean* result);

    LookingAt(
        [out] Boolean* result);

    Matches(
        [out] Boolean* result);

    Pattern(
        [out] IPattern** pattern);

    Region(
        [in] Integer start,
        [in] Integer end);

    RegionStart(
        [out] Integer* start);

    RegionEnd(
        [out] Integer* end);

    ReplaceAll(
        [in] String replacement,
        [out] String* str);

    ReplaceFirst(
        [in] String replacement,
        [out] String* str);

    RequireEnd(
        [out] Boolean* result);

    Reset();

    Reset(
        [in] ICharSequence* input);

    Start(
        [out] Integer* index);

    Start(
        [in] Integer group,
        [out] Integer* index);

    Start(
        [in] String name,
        [out] Integer* index);

    ToMatchResult(
        [out] IMatchResult** result);

    UseAnchoringBounds(
        [in] Boolean value);

    UsePattern(
        [in] IPattern* newPattern);

    UseTransparentBounds(
        [in] Boolean value);
}

[
    uuid(393528c5-7d0a-4304-bd78-c229ebd64a34),
    version(0.1.0)
]
interface IMatcherFactory
{
    QuoteReplacement(
        [in] String s,
        [out] String* str);
}

}
}
}
