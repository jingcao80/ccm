//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {
namespace calendar {

/*
 * @Involve interface ccm::util::calendar::IBaseCalendar
 * @Involve interface ccm::util::calendar::ICalendarSystem
 */
[
    uuid(56b39c04-1748-42e8-901d-64449245f389),
    version(0.1.0)
]
interface ILocalGregorianCalendar
{
    IsLeapYear(
        [in] Integer gregorianYear,
        [out] Boolean* leapYear);

    IsLeapYear(
        [in] IEra* era,
        [in] Integer year,
        [out] Boolean* leapYear);
}

}
}
}
