//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace core {

[
    uuid(21107670-c69c-4bab-b7a2-476469271786),
    version(0.1.0)
]
interface ICharSequence
{
    GetCharAt(
        [in] Integer index,
        [out] Char* c);

    GetLength(
        [out] Integer* number);

    SubSequence(
        [in] Integer start,
        [in] Integer end,
        [out] ICharSequence** subcsq);

    ToString(
        [out] String* str);
}

}
}