//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::core::ICharSequence;

namespace como {
namespace io {

/**
 * @Involve interface como::core::IAppendable;
 * @Involve interface como::io::ICloseable;
 * @Involve interface como::io::IFlushable;
 * @involve interface como::core::IAutoCloseable
 */
[
    uuid(cca035d8-6f23-4eac-a581-294d5ff8c41f),
    version(0.1.0)
]
interface IWriter
{
    Append(
        [in] ICharSequence* csq);

    Append(
        [in] ICharSequence* csq,
        [in] Integer start,
        [in] Integer end);

    Append(
        [in] Char c);

    Close();

    Flush();

    Write(
        [in] Integer c);

    Write(
        [in] Array<Char> buffer);

    Write(
        [in] Array<Char> buffer,
        [in] Integer off,
        [in] Integer len);

    Write(
        [in] String str);

    Write(
        [in] String str,
        [in] Integer off,
        [in] Integer len);
}

}
}
