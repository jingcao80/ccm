//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {

/*
 * @Involve interface ccm::util::ICalendar
 * @Involve interface ccm::io::ISerializable
 * @Involve interface ccm::core::ICloneable
 * @Involve interface ccm::core::IComparable
 */
[
    uuid(7eab4e43-ab92-4309-a542-55d17a8dd6da),
    version(0.1.0)
]
interface IJapaneseImperialCalendar
{
    /**
     * The ERA constant designating the era before Meiji.
     */
    const Integer BEFORE_MEIJI = 0;

    /**
     * The ERA constant designating the Meiji era.
     */
    const Integer MEIJI = 1;

    /**
     * The ERA constant designating the Taisho era.
     */
    const Integer TAISHO = 2;

    /**
     * The ERA constant designating the Showa era.
     */
    const Integer SHOWA = 3;

    /**
     * The ERA constant designating the Heisei era.
     */
    const Integer HEISEI = 4;
}

}
}
