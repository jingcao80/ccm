//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::core::IAppendable;
interface ccm::util::ILocale;

namespace ccm {
namespace util {

/*
 * @Involve interface ccm::io::ICloseable
 * @Involve interface ccm::io::IFlushable
 * @Involve interface ccm::core::IAutoCloseable
 */
[
    uuid(20aae661-0408-4d5e-a0ef-77e433774fac),
    version(0.1.0)
]
interface IFormatter
{
    Close();

    Flush();

    Format(
        [in] String format,
        [in] Array<IInterface*>* args);

    Format(
        [in] ILocale* l,
        [in] String format,
        [in] Array<IInterface*>* args);

    GetIoException(
        [out] ECode* ec);

    GetLocale(
        [out] ILocale** locale);

    GetOut(
        [out] IAppendable** output);

    ToString(
        [out] String* str);
}

}
}
