//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace io {

/*
 * @Involve interface como::io::IBuffer;
 * @Involve interface como::core::IComparable;
 */
[
    uuid(017a5ce6-c447-4245-b1da-fc0d41c4e256),
    version(0.1.0)
]
interface IIntegerBuffer
{
    AsReadOnlyBuffer(
        [out] IIntegerBuffer&& buffer);

    Compact();

    Duplicate(
        [out] IIntegerBuffer&& buffer);

    Get(
        [out] Integer& i);

    Get(
        [in] Integer index,
        [out] Integer& i);

    Get(
        [out] Array<Integer>& dst);

    Get(
        [out] Array<Integer>& dst,
        [in] Integer offset,
        [in] Integer length);

    GetOrder(
        [out] IByteOrder&& bo);

    HasArray(
        [out] Boolean& result);

    Put(
        [in] Integer i);

    Put(
        [in] Integer index,
        [in] Integer i);

    Put(
        [in] Array<Integer> src);

    Put(
        [in] Array<Integer> src,
        [in] Integer offset,
        [in] Integer length);

    Put(
        [in] IIntegerBuffer* src);

    Slice(
        [out] IIntegerBuffer&& buffer);
}

}
}
