//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::util::ILocale;
interface ccm::util::ITimeZone;
interface ccm::util::calendar::ICalendarDate;

namespace ccm {
namespace util {
namespace calendar {

[
    uuid(38c2ed16-4b95-4936-8eab-d418362dd202),
    version(0.1.0)
]
interface IEra
{
    GetAbbreviation(
        [out] String* abbr);

    GetDiaplayAbbreviation(
        [in] ILocale* locale,
        [out] String* abbr);

    GetDisplayName(
        [in] ILocale* locale,
        [out] String* name);

    GetName(
        [out] String* name);

    GetSince(
        [in] ITimeZone* zone,
        [out] Long* time);

    GetSinceDate(
        [out] ICalendarDate** date);

    IsLocalTime(
        [out] Boolean* result);
}

}
}
}
