//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::core::IBoolean;
interface ccm::core::IStringBuffer;
interface ccm::text::IFieldPosition;
interface ccm::text::INumberFormat;
interface ccm::text::IParsePosition;
interface ccm::util::ICalendar;
interface ccm::util::IDate;
interface ccm::util::ILocale;
interface ccm::util::ITimeZone;

namespace ccm {
namespace text {

/*
 * @Involve interface ccm::text::IFormatField
 * @Involve interface ccm::text::IAttributedCharacterIteratorAttribute;
 */
[
    uuid(09b0ec7d-890c-4dda-80dd-e2c32807eda6),
    version(0.1.0)
]
interface IDateFormatField
{
    GetCalendarField(
        [out] Integer* calendarField);
}

/*
 * @Involve interface ccm::text::IFormat;
 * @Involve interface ccm::io::ISerializable;
 * @Involve interface ccm::core::ICloneable;
 */
[
    uuid(4f4122b6-8d1a-4454-ac93-22e858ec23c8),
    version(0.1.0)
]
interface IDateFormat
{
    /**
     * Useful constant for ERA field alignment.
     */
    const Integer ERA_FIELD = 0;

    /**
     * Useful constant for YEAR field alignment.
     */
    const Integer YEAR_FIELD = 1;

    /**
     * Useful constant for MONTH field alignment.
     */
    const Integer MONTH_FIELD = 2;

    /**
     * Useful constant for DATE field alignment.
     */
    const Integer DATE_FIELD = 3;

    /**
     * Useful constant for one-based HOUR_OF_DAY field alignment.
     * HOUR_OF_DAY1_FIELD is used for the one-based 24-hour clock.
     * For example, 23:59 + 01:00 results in 24:59.
     */
    const Integer HOUR_OF_DAY1_FIELD = 4;

    /**
     * Useful constant for zero-based HOUR_OF_DAY field alignment.
     * HOUR_OF_DAY0_FIELD is used for the zero-based 24-hour clock.
     * For example, 23:59 + 01:00 results in 00:59.
     */
    const Integer HOUR_OF_DAY0_FIELD = 5;

    /**
     * Useful constant for MINUTE field alignment.
     */
    const Integer MINUTE_FIELD = 6;

    /**
     * Useful constant for SECOND field alignment.
     */
    const Integer SECOND_FIELD = 7;

    /**
     * Useful constant for MILLISECOND field alignment.
     */
    const Integer MILLISECOND_FIELD = 8;

    /**
     * Useful constant for DAY_OF_WEEK field alignment.
     */
    const Integer DAY_OF_WEEK_FIELD = 9;

    /**
     * Useful constant for DAY_OF_YEAR field alignment.
     */
    const Integer DAY_OF_YEAR_FIELD = 10;

    /**
     * Useful constant for DAY_OF_WEEK_IN_MONTH field alignment.
     */
    const Integer DAY_OF_WEEK_IN_MONTH_FIELD = 11;

    /**
     * Useful constant for WEEK_OF_YEAR field alignment.
     */
    const Integer WEEK_OF_YEAR_FIELD = 12;

    /**
     * Useful constant for WEEK_OF_MONTH field alignment.
     */
    const Integer WEEK_OF_MONTH_FIELD = 13;

    /**
     * Useful constant for AM_PM field alignment.
     */
    const Integer AM_PM_FIELD = 14;

    /**
     * Useful constant for one-based HOUR field alignment.
     * HOUR1_FIELD is used for the one-based 12-hour clock.
     * For example, 11:30 PM + 1 hour results in 12:30 AM.
     */
    const Integer HOUR1_FIELD = 15;

    /**
     * Useful constant for zero-based HOUR field alignment.
     * HOUR0_FIELD is used for the zero-based 12-hour clock.
     * For example, 11:30 PM + 1 hour results in 00:30 AM.
     */
    const Integer HOUR0_FIELD = 16;

    /**
     * Useful constant for TIMEZONE field alignment.
     */
    const Integer TIMEZONE_FIELD = 17;

    /**
     * Constant for full style pattern.
     */
    const Integer FULL = 0;

    /**
     * Constant for long style pattern.
     */
    const Integer LONG = 1;

    /**
     * Constant for medium style pattern.
     */
    const Integer MEDIUM = 2;

    /**
     * Constant for short style pattern.
     */
    const Integer SHORT = 3;

    /**
     * Constant for default style pattern.  Its value is MEDIUM.
     */
    const Integer DEFAULT = MEDIUM;

    Format(
        [in] IDate* date,
        [out] String* result);

    Format(
        [in] IDate* date,
        [in, out] IStringBuffer* toAppendTo,
        [in] IFieldPosition* pos);

    GetCalendar(
        [out] ICalendar** calendar);

    GetNumberFormat(
        [out] INumberFormat** format);

    GetTimeZone(
        [out] ITimeZone** timezone);

    IsLenient(
        [out] Boolean* lenient);

    Parse(
        [in] String source,
        [out] IDate** date);

    Parse(
        [in] String source,
        [in] IParsePosition* pos,
        [out] IDate** date);

    ParseObject(
        [in] String source,
        [in] IParsePosition* pos,
        [out] IInterface** object);

    SetCalendar(
        [in] ICalendar* newCalendar);

    SetLenient(
        [in] Boolean lenient);

    SetNumberFormat(
        [in] INumberFormat* newNumberFormat);

    SetTimeZone(
        [in] ITimeZone* timezone);
}

[
    uuid(70d5b2d6-8ac6-461a-bf2b-dd12826584fc),
    version(0.1.0)
]
interface IDateFormatFactory
{
    GetAvailableLocales(
        [out, callee] Array<ILocale*>* locales);

    GetDateInstance(
        [out] IDateFormat** instance);

    GetDateInstance(
        [in] Integer style,
        [out] IDateFormat** instance);

    GetDateInstance(
        [in] Integer style,
        [in] ILocale* locale,
        [out] IDateFormat** instance);

    GetDateTimeInstance(
        [out] IDateFormat** instance);

    GetDateTimeInstance(
        [in] Integer dateStyle,
        [in] Integer timeStyle,
        [out] IDateFormat** instance);

    GetDateTimeInstance(
        [in] Integer dateStyle,
        [in] Integer timeStyle,
        [in] ILocale* locale,
        [out] IDateFormat** instance);

    GetInstance(
        [out] IDateFormat** instance);

    GetTimeInstance(
        [out] IDateFormat** instance);

    GetTimeInstance(
        [in] Integer style,
        [out] IDateFormat** instance);

    GetTimeInstance(
        [in] Integer style,
        [in] ILocale* locale,
        [out] IDateFormat** instance);

    Set24HourTimePref(
        [in] IBoolean* is24Hour);
}

}
}
