//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::core::INumber;
interface ccm::core::IStringBuffer;
interface ccm::text::IFieldPosition;
interface ccm::text::IParsePosition;

namespace ccm {
namespace text {

/*
 * @Involve interface ccm::text::IFormat;
 * @Involve interface ccm::io::ISerializable;
 * @Involve interface ccm::core::ICloneable;
 */
[
    uuid(69ff7998-7fb1-4f1b-940d-30ad8d233113),
    version(0.1.0)
]
interface INumberFormat
{
    Format(
        [in] Long number,
        [in, out] IStringBuffer* toAppendTo,
        [in] IFieldPosition* pos);

    Format(
        [in] Double number,
        [in, out] IStringBuffer* toAppendTo,
        [in] IFieldPosition* pos);

    Parse(
        [in] String source,
        [out] INumber** number);

    Parse(
        [in] String source,
        [in] IParsePosition* parsePosition,
        [out] INumber** number);

    SetGroupingUsed(
        [in] Boolean value);

    SetMaximumIntegerDigits(
        [in] Integer newValue);

    SetMinimumIntegerDigits(
        [in] Integer newValue);
}

}
}
