//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {

/*
 * @Involve interface ccm::util::IIterator
 */
[
    uuid(e8665718-bf0d-4054-850c-a30098de04b8),
    version(0.1.0)
]
interface IListIterator
{
    Add(
        [in] IInterface* object);

    Next(
        [out] IInterface** object = nullptr);

    GetNextIndex(
        [out] Integer* index);

    Previous(
        [out] IInterface** object = nullptr);

    GetPreviousIndex(
        [out] Integer* index);

    HasNext(
        [out] Boolean* result);

    HasPrevious(
        [out] Boolean* result);

    Remove();

    Set(
        [in] IInterface* object);
}

}
}
