//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::security::IPermission;

namespace como {
namespace core {

[
    uuid(a8d886cf-a4f1-4733-b5ff-a670789b9c25),
    version(0.1.0)
]
interface ISecurityManager
{
    CheckDelete(
        [in] String file);

    CheckExec(
        [in] String file);

    CheckPermission(
        [in] IPermission* perm);

    CheckPropertyAccess(
        [in] String key);

    CheckRead(
        [in] String file);

    CheckWrite(
        [in] String file);
}

}
}
