//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {

/**
 * @Involve interface como::util::IMap
 * @Involve interface como::core::ICloneable
 * @Involve interface como::io::ISerializable
 */
[
    uuid(3b25617c-5ccc-428c-8daf-1bdc855ce1a8),
    version(0.1.0)
]
interface IHashMap
{
    Clear();

    Clone(
        [in] InterfaceID iid,
        [out] IInterface** obj);

    ContainsKey(
        [in] IInterface* key,
        [out] Boolean* result);

    ContainsValue(
        [in] IInterface* value,
        [out] Boolean* result);

    Equals(
        [in] IInterface* obj,
        [out] Boolean& result);

    Get(
        [in] IInterface* key,
        [out] IInterface** value);

    GetEntrySet(
        [out] ISet** entries);

    GetHashCode(
        [out] Integer& hash);

    GetKeySet(
        [out] ISet** keys);

    GetSize(
        [out] Integer* size);

    GetValues(
        [out] ICollection** values);

    IsEmpty(
        [out] Boolean* result);

    Put(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    PutAll(
        [in] IMap* m);

    PutIfAbsent(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    Remove(
        [in] IInterface* key,
        [out] IInterface** prevValue = nullptr);
}

}
}
