//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace core {

[
    uuid(b25cfd17-1013-406e-b0cd-74be7637571c),
    version(0.1.0)
]
interface IThreadGroup
{
    ActiveCount(
        [out] Integer* count);

    ActiveGroupCount(
        [out] Integer* count);

    // @hide
    Add(
        [in] IThread* t);

    // @hide
    AddUnstarted();

    CheckAccess();

    Destroy();

    Enumerate(
        [out] Array<IThread*>& list,
        [out] Integer* count);

    Enumerate(
        [out] Array<IThread*>& list,
        [in] Boolean recurse,
        [out] Integer* count);

    Enumerate(
        [out] Array<IThreadGroup*>& list,
        [out] Integer* count);

    Enumerate(
        [out] Array<IThreadGroup*>& list,
        [in] Boolean recurse,
        [out] Integer* count);

    GetMaxPriority(
        [out] Integer* priority);

    GetName(
        [out] String* name);

    GetParent(
        [out] IThreadGroup** parent);

    Interrupt();

    IsDaemon(
        [out] Boolean* daemon);

    IsDestroyed(
        [out] Boolean* destroyed);

    List();

    ParentOf(
        [in] IThreadGroup* g,
        [out] Boolean* result);

    Resume();

    SetDaemon(
        [in] Boolean daemon);

    SetMaxPriority(
        [in] Integer pri);

    Stop();

    Suspend();

    // @hide
    ThreadStartFailed(
        [in] IThread* t);

    // @hide
    ThreadTerminated(
        [in] IThread* t);
}

}
}
