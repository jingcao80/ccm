//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "como/net/IDatagramPacket.cdl"
include "como/net/IDatagramSocket.cdl"
include "como/net/IInetAddress.cdl"
include "como/net/IInetSocketAddress.cdl"
include "como/net/ISocket.cdl"
include "como/net/ISocketAddress.cdl"
include "como/net/IURI.cdl"
include "como/net/IURL.cdl"
