//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace core {

const Integer E_ILLEGAL_MONITOR_STATE_EXCEPTION = 0x80010100;
const Integer E_INTERRUPTED_EXCEPTION = 0x80010101;
const Integer E_NULL_POINTER_EXCEPTION = 0x80010102;
const Integer E_ILLEGAL_THREAD_STATE_EXCEPTION = 0x80010103;
const Integer E_STRING_INDEX_OUT_OF_BOUNDS_EXCEPTION = 0x80010104;
const Integer E_INDEX_OUT_OF_BOUNDS_EXCEPTION = 0x80010105;
const Integer E_NUMBER_FORMAT_EXCEPTION = 0x80010106;
const Integer E_ILLEGAL_STATE_EXCEPTION = 0x80010107;
const Integer E_ARRAY_INDEX_OUT_OF_BOUNDS_EXCEPTION = 0x80010108;
const Integer E_ARITHMETIC_EXCEPTION = 0x80010109;
const Integer E_CLASS_CAST_EXCEPTION = 0x8001010a;

}
}
