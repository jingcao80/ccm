//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::text::IDateFormatSymbols;
interface como::util::IDate;

namespace como {
namespace text {

/*
 * @Involve interface como::text::IDateFormat;
 * @Involve interface como::text::IFormat;
 * @Involve interface como::io::ISerializable;
 * @Involve interface como::core::ICloneable;
 */
[
    uuid(e2b13317-e567-4a78-96d1-caacffa88817),
    version(0.1.0)
]
interface ISimpleDateFormat
{
    ApplyLocalizedPattern(
        [in] String pattern);

    ApplyPattern(
        [in] String pattern);

    Get2DigitYearStart(
        [out] IDate&& startDate);

    Set2DigitYearStart(
        [in] IDate* startDate);

    SetDateFormatSymbols(
        [in] IDateFormatSymbols* newFormatSymbols);

    ToLocalizedPattern(
        [out] String& pattern);

    ToPattern(
        [out] String& pattern);
}

}
}
