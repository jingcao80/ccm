//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {

interface IIterator;

[
    uuid(2618a380-071b-440b-84b7-d3ac4a3de3ad),
    version(0.1.0)
]
interface ICollection
{
    Add(
        [in] IInterface* obj,
        [out] Boolean* changed = nullptr);

    AddAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    Clear();

    Contains(
        [in] IInterface* obj,
        [out] Boolean* result);

    ContainsAll(
        [in] ICollection* c,
        [out] Boolean* result);

    Equals(
        [in] IInterface* obj,
        [out] Boolean* result);

    GetHashCode(
        [out] Integer* hash);

    GetIterator(
        [out] IIterator** it);

    GetSize(
        [out] Integer* size);

    IsEmpty(
        [out] Boolean* empty);

    Remove(
        [in] IInterface* obj,
        [out] Boolean* changed = nullptr);

    RemoveAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    RetainAll(
        [in] ICollection* c,
        [out] Boolean* changed = nullptr);

    ToArray(
        [in] InterfaceID iid,
        [out, callee] Array<IInterface*>* objs);
}

}
}
