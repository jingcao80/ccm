//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

[
    uuid(3657416d-4638-4843-a0b9-eb7ef1794495),
    uri("http://como.org/component/library/libcore.so")
]
module libcore
{

include "como/core.cdl"
include "como/io.cdl"
include "como/core2.cdl"
include "como/math.cdl"
include "como/misc.cdl"
include "como/net.cdl"
include "como/security.cdl"
include "como/core3.cdl"
include "como/text.cdl"
include "como/util.cdl"
include "comort/system.cdl"
include "libcore/icu.cdl"
include "libcore/io.cdl"
include "libcore/util.cdl"
include "pisces/icu.cdl"
include "pisces/system.cdl"

}
