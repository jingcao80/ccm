//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::math::IBigInteger;
interface como::math::IMathContext;
enum como::math::RoundingMode;

namespace como {
namespace math {

[
    uuid(51317f66-2236-494c-9eef-da37c95a2845),
    version(0.1.0)
]
interface IBigDecimal
{
    const Integer ROUND_UP = 0;

    const Integer ROUND_DOWN = 1;

    const Integer ROUND_CEILING = 2;

    const Integer ROUND_FLOOR = 3;

    const Integer ROUND_HALF_UP = 4;

    const Integer ROUND_HALF_DOWN = 5;

    const Integer ROUND_HALF_EVEN = 6;

    const Integer ROUND_UNNECESSARY = 7;

    Abs(
        [out] IBigDecimal&& value);

    Abs(
        [in] IMathContext* mc,
        [out] IBigDecimal&& value);

    Add(
        [in] IBigDecimal* augend,
        [out] IBigDecimal&& result);

    Add(
        [in] IBigDecimal* augend,
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    ByteValueExact(
        [out] Byte& value);

    Divide(
        [in] IBigDecimal* divisor,
        [out] IBigDecimal&& result);

    Divide(
        [in] IBigDecimal* divisor,
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    Divide(
        [in] IBigDecimal* divisor,
        [in] Integer roundingMode,
        [out] IBigDecimal&& result);

    Divide(
        [in] IBigDecimal* divisor,
        [in] RoundingMode roundingMode,
        [out] IBigDecimal&& result);

    Divide(
        [in] IBigDecimal* divisor,
        [in] Integer scale,
        [in] Integer roundingMode,
        [out] IBigDecimal&& result);

    Divide(
        [in] IBigDecimal* divisor,
        [in] Integer scale,
        [in] RoundingMode roundingMode,
        [out] IBigDecimal&& result);

    DivideAndRemainder(
        [in] IBigDecimal* divisor,
        [out, callee] Array<IBigDecimal*>* quotAndRem);

    DivideAndRemainder(
        [in] IBigDecimal* divisor,
        [in] IMathContext* mc,
        [out, callee] Array<IBigDecimal*>* quotAndRem);

    DivideToIntegralValue(
        [in] IBigDecimal* divisor,
        [out] IBigDecimal&& result);

    DivideToIntegralValue(
        [in] IBigDecimal* divisor,
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    IntegerValueExact(
        [out] Integer& value);

    LongValueExact(
        [out] Long& value);

    Max(
        [in] IBigDecimal* value,
        [out] IBigDecimal&& result);

    Min(
        [in] IBigDecimal* value,
        [out] IBigDecimal&& result);

    MovePointLeft(
        [in] Integer n,
        [out] IBigDecimal&& value);

    MovePointRight(
        [in] Integer n,
        [out] IBigDecimal&& value);

    Multiply(
        [in] IBigDecimal* multiplicand,
        [out] IBigDecimal&& result);

    Multiply(
        [in] IBigDecimal* multiplicand,
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    Negate(
        [out] IBigDecimal&& value);

    Negate(
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    Plus(
        [out] IBigDecimal&& value);

    Plus(
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    Pow(
        [in] Integer n,
        [out] IBigDecimal&& value);

    Pow(
        [in] Integer n,
        [in] IMathContext* mc,
        [out] IBigDecimal&& value);

    Precision(
        [out] Integer& precision);

    Remainder(
        [in] IBigDecimal* divisor,
        [out] IBigDecimal&& result);

    Remainder(
        [in] IBigDecimal* divisor,
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    Round(
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    Scale(
        [out] Integer& scale);

    ScaleByPowerOfTen(
        [in] Integer n,
        [out] IBigDecimal&& value);

    SetScale(
        [in] Integer newScale,
        [out] IBigDecimal&& value);

    SetScale(
        [in] Integer newScale,
        [in] Integer roundingMode,
        [out] IBigDecimal&& result);

    SetScale(
        [in] Integer newScale,
        [in] RoundingMode roundingMode,
        [out] IBigDecimal&& result);

    ShortValueExact(
        [out] Short& value);

    Signum(
        [out] Integer& sign);

    StripTrailingZeros(
        [out] IBigDecimal&& value);

    Subtract(
        [in] IBigDecimal* subtrahend,
        [out] IBigDecimal&& result);

    Subtract(
        [in] IBigDecimal* subtrahend,
        [in] IMathContext* mc,
        [out] IBigDecimal&& result);

    ToBigInteger(
        [out] IBigInteger&& value);

    ToBigIntegerExact(
        [out] IBigInteger&& value);

    ToEngineeringString(
        [out] String& desc);

    ToPlainString(
        [out] String& desc);

    Ulp(
        [out] IBigDecimal&& value);

    UnscaledValue(
        [out] IBigInteger&& value);
}

}
}
