//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "libcore/util/IBasicLruCache.cdl"
include "libcore/util/IZoneInfo.cdl"
include "libcore/util/IZoneInfoDB.cdl"

namespace libcore {
namespace util {

[
    uuid(b9bc96e1-babc-46c0-86f4-79c914e06ef9),
    version(0.1.0)
]
coclass CZoneInfoWallTime
{
    Constructor();

    interface IZoneInfoWallTime;
}

}
}
