//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

[
    uuid(3a58f162-2708-4f66-bd21-faaef914063b),
    uri("http://ccm.org/component/test/NestedInterfaceTest.so")
]
module NestedInterfaceTest
{

namespace ccm {
namespace test {

[
    uuid(d7542341-9da2-4288-bca5-50cfebfe6700),
    version(0.1.0)
]
interface IFooBar
{
    [
        uuid(19cfe29d-55cd-4572-a1b0-9167103aff28),
        version(0.1.0)
    ]
    interface IFoo
    {
        Foo1();

        Foo2();
    }

    FooBar1();

    FooBar2();

    [
        uuid(9b408e72-2787-4465-b03a-5ccbaf4cd2b8),
        version(0.1.0)
    ]
    interface IBar
    {
        Bar1();

        Bar2(
            [in] IFoo* foo);
    }

    FooBar3();
}

[
    uuid(9050982a-7f29-4630-922f-55be9e6d437e),
    version(0.1.0)
]
coclass CFooBar
{
    Constructor(
        [in] IFooBar::IFoo* foo);

    interface IFooBar::IFoo;
    interface IFooBar::IBar;
}

}
}

}
