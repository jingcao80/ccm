//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ccm/text/Exceptions.cdl"
include "ccm/text/IAttributedCharacterIterator.cdl"
include "ccm/text/IAttributedString.cdl"
include "ccm/text/ICharacterIterator.cdl"
include "ccm/text/IDateFormat.cdl"
include "ccm/text/IDateFormatSymbols.cdl"
include "ccm/text/IDecimalFormat.cdl"
include "ccm/text/IDecimalFormatSymbols.cdl"
include "ccm/text/IFieldPosition.cdl"
include "ccm/text/IFormat.cdl"
include "ccm/text/INumberFormat.cdl"
include "ccm/text/IParsePosition.cdl"
include "ccm/text/ISimpleDateFormat.cdl"

interface ccm::core::ICloneable;
interface ccm::io::ISerializable;
interface ccm::util::ILocale;
interface ccm::util::IMap;

namespace ccm {
namespace text {

[
    uuid(812928e8-cbef-4bbe-a33d-792341c3d681),
    version(0.1.0)
]
coclass CAttributedCharacterIteratorAttribute
{
    Constructor() = delete;

    interface IAttributedCharacterIteratorAttribute;
    interface ISerializable;
}

[
    uuid(d90f0463-63bb-43dd-8ae6-69152b0fcbd1),
    version(0.1.0)
]
coclass CAttributedString
{
    Constructor(
        [in] Array<IAttributedCharacterIterator*> iterators);

    Constructor(
        [in] String text);

    Constructor(
        [in] String text,
        [in] IMap* attributes);

    Constructor(
        [in] IAttributedCharacterIterator* text);

    Constructor(
        [in] IAttributedCharacterIterator* text,
        [in] Integer beginIndex,
        [in] Integer endIndex);

    Constructor(
        [in] IAttributedCharacterIterator* text,
        [in] Integer beginIndex,
        [in] Integer endIndex,
        [in] Array<IAttributedCharacterIteratorAttribute*> attributes);

    interface IAttributedString;
}

[
    uuid(43ac1b62-c9d8-4345-a293-f27cf49427f0),
    version(0.1.0)
]
coclass CDateFormatField
{
    Constructor() = delete;

    interface IDateFormatField;
    interface IFormatField;
    interface IAttributedCharacterIteratorAttribute;
    interface ISerializable;
}

[
    uuid(5eade1e5-5963-4f1b-bfc1-9f1f9ae4b52f),
    version(0.1.0)
]
coclass CDecimalFormat
{
    Constructor();

    Constructor(
        [in] String pattern);

    Constructor(
        [in] String pattern,
        [in] IDecimalFormatSymbols* symbols);

    interface ccm::text::IDecimalFormat;
    interface ccm::text::INumberFormat;
    interface ccm::text::IFormat;
    interface ccm::io::ISerializable;
    interface ccm::core::ICloneable;
}

[
    uuid(81e790a2-a790-4776-b726-8502d7271000),
    version(0.1.0)
]
coclass CDecimalFormatSymbols
{
    Constructor();

    Constructor(
        [in] ILocale* locale);

    interface IDecimalFormatSymbols;
    interface ICloneable;
    interface ISerializable;
}

[
    uuid(6081b56d-7a1b-4676-8122-f28f2e319c49),
    version(0.1.0)
]
coclass CFieldPosition
{
    Constructor(
        [in] Integer field);

    Constructor(
        [in] IFormatField* attribute);

    Constructor(
        [in] IFormatField* attribute,
        [in] Integer field);

    interface IFieldPosition;
}

[
    uuid(cc8abe8d-754f-4020-8c93-fbcb73887861),
    version(0.1.0)
]
coclass CNumberFormatFactory
{
    interface INumberFormatFactory;
}

[
    uuid(5dd60879-0252-4319-a926-70517a5484e1),
    version(0.1.0)
]
coclass CParsePosition
{
    Constructor(
        [in] Integer index);

    interface IParsePosition;
}

[
    uuid(abcdea41-9127-42d0-a5e0-ac4f1bb9d249),
    version(0.1.0)
]
coclass CSimpleDateFormat
{
    Constructor();

    Constructor(
        [in] String pattern);

    Constructor(
        [in] String pattern,
        [in] ILocale* locale);

    Constructor(
        [in] String pattern,
        [in] IDateFormatSymbols* formatSymbols);

    interface ISimpleDateFormat;
    interface IDateFormat;
    interface IFormat;
    interface ISerializable;
    interface ICloneable;
}

}
}
