//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace util {

[
    uuid(c548a9de-f3d8-4acb-83f3-00c65c1b56b2),
    version(0.1.0)
]
interface IComparator
{
    Compare(
        [in] IInterface* o1,
        [in] IInterface* o2,
        [out] Integer* result);

    Equals(
        [in] IInterface* obj,
        [out] Boolean* isEqual);
}

}
}
