//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {

/*
 * @Involve interface como::io:ISerializable
 */
[
    uuid(b262d480-e46b-49c2-acba-98478d810a12),
    version(0.1.0)
]
interface IRandom
{
    NextBoolean(
        [out] Boolean& value);

    NextBytes(
        [out] Array<Byte>& bytes);

    NextDouble(
        [out] Double& value);

    NextFloat(
        [out] Float& value);

    NextGaussian(
        [out] Double& value);

    NextInteger(
        [out] Integer& value);

    NextInteger(
        [in] Integer bound,
        [out] Integer& value);

    NextLong(
        [out] Long& value);

    SetSeed(
        [in] Long seed);
}

}
}
