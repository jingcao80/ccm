//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

/**
 * Test parsing module.
 */

[
    uuid(6c69c8bc-b62d-4dad-811b-26f73cd2aaa7),
    url("http://ccm.org/components/test/test_module.so"),
    description("This is the definition of module TestModule.")
]
module TestModule
{

include "interfaceTests.cdl"
include "coclassTests.cdl"

}
