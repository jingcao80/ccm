//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {
namespace regex {

[
    uuid(37d33b90-45d9-4b01-88e8-982e7e830c21),
    version(0.1.0)
]
interface IMatchResult
{
    End(
        [out] Integer& index);

    End(
        [in] Integer group,
        [out] Integer& index);

    Group(
        [out] String& subseq);

    Group(
        [in] Integer group,
        [out] String& subseq);

    GroupCount(
        [out] Integer& number);

    Start(
        [out] Integer& index);

    Start(
        [in] Integer group,
        [out] Integer& index);
}

}
}
}
