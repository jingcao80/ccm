//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::util::ISet;

namespace ccm {
namespace util {

[
    uuid(b77f3ad5-3301-486b-a529-24fe27caa151),
    version(0.1.0)
]
interface ILocaleCategory
{
    GetLanguageKey(
        [out] String* key);

    GetScriptKey(
        [out] String* key);

    GetCountryKey(
        [out] String* key);

    GetVariantKey(
        [out] String* key);
}

/*
 * @Involve ccm::core::ICloneable
 * @Involve ccm::io::ISerializable
 */
[
    uuid(e23a921a-6d45-4b08-89e3-f09778118022),
    version(0.1.0)
]
interface ILocale
{
    GetCountry(
        [out] String* country);

    GetExtension(
        [in] Char key,
        [out] String* extension);

    GetExtensionKeys(
        [out] ISet** keys);

    GetLanguage(
        [out] String* language);

    GetScript(
        [out] String* script);

    GetUnicodeLocaleAttributes(
        [out] ISet** attrs);

    GetUnicodeLocaleKeys(
        [out] ISet** keys);

    GetUnicodeLocaleType(
        [in] String key,
        [out] String* type);

    GetVariant(
        [out] String* variant);

    ToLanguageTag(
        [out] String* langTag);
}

}
}
