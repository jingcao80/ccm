//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace util {
namespace concurrent {
namespace atomic {

/*
 * @Involve interface como::io::ISerializable
 */
[
    uuid(2251febf-a611-4962-9d23-b6e505a3d4d8),
    version(0.1.0)
]
interface IAtomicBoolean
{
    CompareAndSet(
        [in] Boolean expect,
        [in] Boolean update,
        [out] Boolean* succeeded = nullptr);

    Get(
        [out] Boolean* value);

    GetAndSet(
        [in] Boolean newValue,
        [out] Boolean* prevValue);

    LzaySet(
        [in] Boolean value);

    Set(
        [in] Boolean value);

    WeakCompareAndSet(
        [in] Boolean expect,
        [in] Boolean update,
        [out] Boolean* succeeded = nullptr);
}

}
}
}
}
