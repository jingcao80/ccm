//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::io::ISerializable;
interface como::security::IGuard;
interface como::security::IPermission;

namespace como {
namespace core {

[
    uuid(106e254e-0909-4238-8db4-2e343715c9ad),
    version(0.1.0)
]
coclass CRuntimePermission
{
    Constructor(
        [in] String name);

    Constructor(
        [in] String name,
        [in] String actions);

    interface IPermission;
    interface IGuard;
    interface ISerializable;
}

}
}
