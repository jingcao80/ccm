//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::security::IPermission;
interface como::util::IEnumeration;

namespace como {
namespace security {

/*
 * @Involve interface como::io::ISerializable
 */
[
    uuid(8bdc918c-d6b9-457b-8d4c-24cdb0a4ed42),
    version(0.1.0)
]
interface IPermissionCollection
{
    Add(
        [in] IPermission* permission);

    GetElements(
        [out] IEnumeration&& elements);

    Implies(
        [in] IPermission* permission,
        [out] Boolean& result);

    IsReadOnly(
        [out] Boolean& readonly);

    SetReadOnly();
}

}
}
