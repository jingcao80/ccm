//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::core::IInteger;

namespace libcore {
namespace icu {

[
    uuid(b3ead832-20d3-43cd-9246-7654f4626ae4),
    version(0.1.0)
]
interface ILocaleData
{
    GetCurrencySymbol(
        [out] String* currencySymbol);

    GetDateFormat(
        [in] Integer style,
        [out] String* dateFormat);

    GetDecimalSeparator(
        [out] Char* decSeparator);

    GetExponentSeparator(
        [out] String* expSeparator);

    GetGroupingSeparator(
        [out] Char* grpSeparator);

    GetFirstDayOfWeek(
        [out] IInteger** day);

    GetInfinity(
        [out] String* infinity);

    GetInternationalCurrencySymbol(
        [out] String* intlCurrencySymbol);

    GetMinimalDaysInFirstWeek(
        [out] IInteger** days);

    GetMinusSign(
        [out] String* sign);

    GetNaN(
        [out] String* nan);

    GetPatternSeparator(
        [out] Char* patSeparator);

    GetPercent(
        [out] String* percent);

    GetPerMill(
        [out] Char* perMill);

    GetTimeFormat(
        [in] Integer style,
        [out] String* timeFormat);

    GetZeroDigit(
        [out] Char* zeroDigit);
}

}
}
