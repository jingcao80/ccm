//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::core::ICharSequence;

namespace como {
namespace util {
namespace regex {

interface IMatcher;

[
    uuid(89258176-0af5-40ce-80bb-0b661dde40bf),
    version(0.1.0)
]
interface IPattern
{
    const Integer UNIX_LINES = 0x01;

    const Integer CASE_INSENSITIVE = 0x02;

    const Integer COMMENTS = 0x04;

    const Integer MULTILINE = 0x08;

    const Integer LITERAL = 0x10;

    const Integer DOTALL = 0x20;

    const Integer UNICODE_CASE = 0x40;

    const Integer CANON_EQ = 0x80;

    Flags(
        [out] Integer& flags);

    Matcher(
        [in] ICharSequence* input,
        [out] IMatcher&& matcher);

    GetPattern(
        [out] String& pattStr);

    Split(
        [in] ICharSequence* input,
        [in] Integer limit,
        [out, callee] Array<String>* strArray);

    Split(
        [in] ICharSequence* input,
        [out, callee] Array<String>* strArray);

    ToString(
        [out] String& pattStr);
}

}
}
}
