//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::util::IEnumeration;

namespace como {
namespace util {
namespace concurrent {

/*
 * @Involve interface como::util::concurrent::IConcurrentMap
 * @Involve interface como::util::IMap
 * @Involve interface como::io::ISerializable
 */
[
    uuid(7f68ef50-b944-403d-a1d3-1fe5c81c094e),
    version(0.1.0)
]
interface IConcurrentHashMap
{
    Clear();

    Contains(
        [in] IInterface* value,
        [out] Boolean* result);

    ContainsKey(
        [in] IInterface* key,
        [out] Boolean* result);

    ContainsValue(
        [in] IInterface* value,
        [out] Boolean* result);

    Elements(
        [out] IEnumeration** elements);

    Equals(
        [in] IInterface* obj,
        [out] Boolean* result);

    Get(
        [in] IInterface* key,
        [out] IInterface** value);

    GetEntrySet(
        [out] ISet** entries);

    GetHashCode(
        [out] Integer* hash);

    GetKeySet(
        [out] ISet** keys);

    GetKeySet(
        [in] IInterface* mappedValue,
        [out] ISet** keys);

    GetMappingCount(
        [out] Long* count);

    GetSize(
        [out] Integer* size);

    GetValues(
        [out] ICollection** values);

    IsEmpty(
        [out] Boolean* result);

    Keys(
        [out] IEnumeration** keys);

    Put(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    PutAll(
        [in] IMap* m);

    PutIfAbsent(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    Remove(
        [in] IInterface* key,
        [out] IInterface** prevValue = nullptr);

    Remove(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] Boolean* result = nullptr);

    Replace(
        [in] IInterface* key,
        [in] IInterface* value,
        [out] IInterface** prevValue = nullptr);

    Replace(
        [in] IInterface* key,
        [in] IInterface* oldValue,
        [in] IInterface* newValue,
        [out] Boolean* result = nullptr);
}

}
}
}
