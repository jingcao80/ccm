//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

/**
 * This file contains the definition of interface ICelestialBody.
 * ICelestialBody stands for all the celestial body in the Universe.
 */

enum CelestialBodyKind
{
    meteor,
    planet,
    satellite,
    star
}

[
    uuid(38fe0857-a480-4d3b-9f6b-1701a760266d),
    version(0.1.0),
    description("This is the definition of ICelestialBody.")
]
interface ICelestialBody
{
    GetName(
        [out] String* name);

    GetKind(
        [out] CelestialBodyKind* kind);

    GetSpace(
        [out] String* universe);

    GetPosition(
        [out] Float* latitude,
        [out] Float* longitude);

    GetSize(
        [out] Double* size);

    GetWeight(
        [out] Double* weight);

    GetAge(
        [out] Integer* age);
}
