//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::security::IPermissionCollection;

namespace como {
namespace security {

/*
 * @Involve interface como::security::IGuard
 * @Involve interface como::io::ISerializable
 */
[
    uuid(93cc3a78-0afc-4b41-999c-aaa643c6e1a3),
    version(0.1.0)
]
interface IPermission
{
    CheckGuard(
        [in] IInterface* object);

    GetActions(
        [out] String* actions);

    GetName(
        [out] String* name);

    Implies(
        [in] IPermission* permission,
        [out] Boolean* result);

    NewPermissionCollection(
        [out] IPermissionCollection** permissions);
}

}
}
