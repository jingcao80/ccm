//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace ccm {
namespace text {

/*
 * @Involve interface ccm::text::INumberFormat;
 * @Involve interface ccm::text::IFormat;
 * @Involve interface ccm::io::ISerializable;
 * @Involve interface ccm::core::ICloneable;
 */
[
    uuid(54f82f1f-4aaf-45b6-891d-77083bff1058),
    version(0.1.0)
]
interface IChoiceFormat
{
    ToPattern(
        [out] String* pattern);
}

}
}
