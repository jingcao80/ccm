//=========================================================================
// Copyright (C) 2018 The C++ Component Model(CCM) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface ccm::util::ISet;

namespace ccm {
namespace util {

[
    uuid(b77f3ad5-3301-486b-a529-24fe27caa151),
    version(0.1.0)
]
interface ILocaleCategory
{
    GetLanguageKey(
        [out] String* key);

    GetScriptKey(
        [out] String* key);

    GetCountryKey(
        [out] String* key);

    GetVariantKey(
        [out] String* key);
}

interface ILocale;

[
    uuid(533f5611-bdc2-4c2a-a6f7-07a9267080c2),
    version(0.1.0)
]
interface ILocaleBuilder
{
    AddUnicodeLocaleAttribute(
        [in] String attribute);

    Build(
        [out] ILocale** locale);

    Clear();

    ClearExtensions();

    RemoveUnicodeLocaleAttribute(
        [in] String attribute);

    SetExtension(
        [in] Char key,
        [in] String value);

    SetLanguage(
        [in] String language);

    SetLanguageTag(
        [in] String languageTag);

    SetLocale(
        [in] ILocale* locale);

    SetRegion(
        [in] String region);

    SetScript(
        [in] String script);

    SetUnicodeLocaleKeyword(
        [in] String key,
        [in] String type);

    SetVariant(
        [in] String variant);
}

/*
 * @Involve ccm::core::ICloneable
 * @Involve ccm::io::ISerializable
 */
[
    uuid(e23a921a-6d45-4b08-89e3-f09778118022),
    version(0.1.0)
]
interface ILocale
{
    GetCountry(
        [out] String* country);

    GetDisplayCountry(
        [out] String* country);

    GetDisplayCountry(
        [in] ILocale* locale,
        [out] String* country);

    GetDisplayLanguage(
        [out] String* language);

    GetDisplayLanguage(
        [in] ILocale* locale,
        [out] String* language);

    GetDisplayName(
        [out] String* name);

    GetDisplayName(
        [in] ILocale* locale,
        [out] String* name);

    GetDisplayScript(
        [out] String* script);

    GetDisplayScript(
        [in] ILocale* inLocale,
        [out] String* script);

    GetDisplayVariant(
        [out] String* variant);

    GetDisplayVariant(
        [in] ILocale* inLocale,
        [out] String* variant);

    GetExtension(
        [in] Char key,
        [out] String* extension);

    GetExtensionKeys(
        [out] ISet** keys);

    GetISO3Country(
        [out] String* country);

    GetISO3Language(
        [out] String* language);

    GetLanguage(
        [out] String* language);

    GetScript(
        [out] String* script);

    GetUnicodeLocaleAttributes(
        [out] ISet** attrs);

    GetUnicodeLocaleKeys(
        [out] ISet** keys);

    GetUnicodeLocaleType(
        [in] String key,
        [out] String* type);

    GetVariant(
        [out] String* variant);

    ToLanguageTag(
        [out] String* langTag);
}

[
    uuid(e7ebb9fa-52aa-470d-bdd6-873bf2c1e87d),
    version(0.1.0)
]
interface ILocaleFactory
{
    GetDefault(
        [out] ILocale** l);
}

}
}
